magic
tech scmos
timestamp 1701546693
<< nwell >>
rect 863 1568 909 1587
rect 923 1584 984 1601
rect 647 1505 731 1506
rect 647 1486 798 1505
rect 809 1487 855 1506
rect 647 1476 752 1486
rect 666 1302 776 1303
rect 855 1302 954 1303
rect 620 1283 776 1302
rect 809 1283 954 1302
rect 967 1283 1013 1302
rect 674 1274 776 1283
rect 855 1274 954 1283
rect 1020 1270 1097 1302
rect 297 1266 361 1267
rect 186 1247 232 1266
rect 257 1247 361 1266
rect 1125 1265 1171 1284
rect 1185 1281 1246 1298
rect 1853 1255 1913 1272
rect 308 1240 361 1247
rect 309 1239 361 1240
rect 1927 1239 1973 1258
rect 1988 1255 2049 1272
rect 2063 1239 2109 1258
rect 2134 1257 2195 1274
rect 2209 1241 2255 1260
rect 2282 1257 2342 1274
rect 2356 1241 2402 1260
rect 2493 1256 2554 1273
rect 2568 1240 2614 1259
rect 2629 1256 2690 1273
rect 2704 1240 2750 1259
rect 2775 1258 2836 1275
rect 2850 1242 2896 1261
rect 2922 1258 2983 1275
rect 2997 1242 3043 1261
rect 376 1200 443 1228
rect 458 1204 504 1223
rect 1852 1147 1913 1164
rect 1927 1131 1973 1150
rect 1996 1147 2057 1164
rect 2071 1131 2117 1150
rect 2145 1149 2206 1166
rect 2220 1133 2266 1152
rect 2290 1150 2351 1167
rect 2365 1134 2411 1153
rect 1545 1077 1606 1094
rect 1618 1062 1664 1081
rect 294 1044 358 1045
rect 183 1025 229 1044
rect 254 1025 358 1044
rect 305 1018 358 1025
rect 678 1019 724 1038
rect 738 1035 799 1052
rect 825 1019 871 1038
rect 885 1035 946 1052
rect 306 1017 358 1018
rect 971 1017 1017 1036
rect 1031 1033 1092 1050
rect 1107 1017 1153 1036
rect 1167 1033 1228 1050
rect 380 1006 403 1011
rect 373 978 440 1006
rect 455 982 501 1001
rect 1544 959 1605 976
rect 2253 967 2314 984
rect 669 912 715 931
rect 729 928 790 945
rect 814 911 860 930
rect 874 927 935 944
rect 1617 943 1663 962
rect 2328 951 2374 970
rect 2389 967 2450 984
rect 2464 951 2510 970
rect 2535 969 2596 986
rect 2610 953 2656 972
rect 2682 969 2743 986
rect 2757 953 2803 972
rect 963 909 1009 928
rect 1023 925 1084 942
rect 1107 909 1153 928
rect 1167 925 1228 942
rect 1390 923 1474 942
rect 2055 908 2101 909
rect 1990 890 2101 908
rect 1990 888 2055 890
rect 49 871 147 872
rect 3 852 147 871
rect 297 859 361 860
rect 49 843 147 852
rect 161 840 232 859
rect 257 840 361 859
rect 1543 855 1604 872
rect 2253 859 2314 876
rect 308 833 361 840
rect 1618 839 1664 858
rect 2328 843 2374 862
rect 2397 859 2458 876
rect 2472 843 2518 862
rect 2546 861 2607 878
rect 2621 845 2667 864
rect 2691 862 2752 879
rect 2766 846 2812 865
rect 309 832 361 833
rect 388 824 406 826
rect 383 821 406 824
rect 376 793 443 821
rect 458 797 504 816
rect 1543 759 1604 776
rect 1616 743 1663 762
rect 297 684 361 685
rect 186 665 232 684
rect 257 665 361 684
rect 308 658 361 665
rect 309 657 361 658
rect 2053 654 2117 655
rect 379 646 406 651
rect 376 618 443 646
rect 458 622 504 641
rect 2009 635 2117 654
rect 2064 628 2117 635
rect 2065 627 2117 628
rect 2139 616 2162 621
rect 2132 588 2199 616
rect 2214 592 2260 611
rect 1461 529 1507 548
rect 1514 519 1598 549
rect 2047 471 2111 472
rect 2003 452 2111 471
rect 2058 445 2111 452
rect 2059 444 2111 445
rect 2133 433 2156 438
rect 1287 396 1333 415
rect 1347 412 1408 429
rect 1433 394 1479 413
rect 1493 410 1554 427
rect 1569 394 1615 413
rect 1629 410 1690 427
rect 2126 405 2193 433
rect 2208 409 2254 428
rect 2035 299 2099 300
rect 1378 282 1451 283
rect 1485 282 1497 284
rect 1716 282 1784 283
rect 1378 263 1500 282
rect 1716 263 1838 282
rect 1991 280 2099 299
rect 2046 273 2099 280
rect 2047 272 2099 273
rect 1378 256 1431 263
rect 1716 256 1769 263
rect 2121 261 2144 266
rect 1378 255 1430 256
rect 1716 255 1768 256
rect 1333 245 1353 249
rect 1333 244 1363 245
rect 1671 244 1694 249
rect 1235 220 1281 239
rect 1296 216 1363 244
rect 1573 220 1619 239
rect 1634 216 1701 244
rect 2114 233 2181 261
rect 2196 237 2242 256
rect 2026 115 2090 116
rect 1982 96 2090 115
rect 2037 89 2090 96
rect 2038 88 2090 89
rect 2112 77 2135 82
rect 2105 49 2172 77
rect 2187 53 2233 72
rect 1429 8 1475 27
rect 1482 -2 1566 28
rect 1255 -125 1301 -106
rect 1315 -109 1376 -92
rect 1401 -127 1447 -108
rect 1461 -111 1522 -94
rect 1537 -127 1583 -108
rect 1597 -111 1658 -94
rect 1346 -239 1419 -238
rect 1453 -239 1465 -237
rect 1684 -239 1752 -238
rect 1346 -258 1468 -239
rect 1684 -258 1806 -239
rect 1346 -265 1399 -258
rect 1684 -265 1737 -258
rect 1346 -266 1398 -265
rect 1684 -266 1736 -265
rect 1301 -277 1330 -272
rect 1639 -277 1668 -272
rect 1203 -301 1249 -282
rect 1264 -305 1331 -277
rect 1541 -301 1587 -282
rect 1602 -305 1669 -277
rect 1429 -443 1475 -424
rect 1482 -453 1566 -423
rect 1255 -576 1301 -557
rect 1315 -560 1376 -543
rect 1401 -578 1447 -559
rect 1461 -562 1522 -545
rect 1537 -578 1583 -559
rect 1597 -562 1658 -545
rect 1346 -690 1419 -689
rect 1453 -690 1465 -688
rect 1684 -690 1752 -689
rect 1346 -709 1468 -690
rect 1684 -709 1806 -690
rect 1346 -716 1399 -709
rect 1684 -716 1737 -709
rect 1346 -717 1398 -716
rect 1684 -717 1736 -716
rect 1301 -728 1330 -723
rect 1639 -727 1668 -723
rect 1639 -728 1669 -727
rect 1203 -752 1249 -733
rect 1264 -756 1331 -728
rect 1541 -752 1587 -733
rect 1602 -756 1669 -728
rect 1420 -893 1466 -874
rect 1473 -903 1557 -873
rect 1246 -1026 1292 -1007
rect 1306 -1010 1367 -993
rect 1392 -1028 1438 -1009
rect 1452 -1012 1513 -995
rect 1528 -1028 1574 -1009
rect 1588 -1012 1649 -995
rect 1337 -1140 1410 -1139
rect 1444 -1140 1456 -1138
rect 1675 -1140 1743 -1139
rect 1337 -1159 1459 -1140
rect 1675 -1159 1797 -1140
rect 1337 -1166 1390 -1159
rect 1675 -1166 1728 -1159
rect 1337 -1167 1389 -1166
rect 1675 -1167 1727 -1166
rect 1292 -1178 1321 -1173
rect 1630 -1178 1653 -1173
rect 1194 -1202 1240 -1183
rect 1255 -1187 1321 -1178
rect 1255 -1206 1322 -1187
rect 1532 -1202 1578 -1183
rect 1593 -1206 1660 -1178
<< ntransistor >>
rect 936 1561 941 1566
rect 959 1561 964 1566
rect 878 1553 883 1558
rect 778 1471 783 1476
rect 835 1472 840 1477
rect 669 1453 674 1458
rect 685 1453 690 1458
rect 701 1453 706 1458
rect 717 1453 722 1458
rect 635 1268 640 1273
rect 824 1268 829 1273
rect 982 1268 987 1273
rect 406 1250 411 1255
rect 424 1250 429 1255
rect 690 1252 695 1257
rect 706 1252 711 1257
rect 722 1252 727 1257
rect 738 1252 743 1257
rect 754 1252 759 1257
rect 883 1252 888 1257
rect 899 1252 904 1257
rect 915 1252 920 1257
rect 931 1252 936 1257
rect 212 1232 217 1237
rect 272 1232 277 1237
rect 1045 1251 1050 1256
rect 1061 1251 1066 1256
rect 1077 1251 1082 1256
rect 1198 1258 1203 1263
rect 1221 1258 1226 1263
rect 1140 1250 1145 1255
rect 1872 1232 1877 1237
rect 1895 1232 1900 1237
rect 323 1211 328 1216
rect 341 1211 346 1216
rect 2008 1232 2013 1237
rect 2031 1232 2036 1237
rect 2154 1234 2159 1239
rect 2177 1234 2182 1239
rect 1953 1224 1958 1229
rect 2089 1224 2094 1229
rect 2301 1234 2306 1239
rect 2324 1234 2329 1239
rect 2235 1226 2240 1231
rect 2513 1233 2518 1238
rect 2536 1233 2541 1238
rect 2382 1226 2387 1231
rect 2649 1233 2654 1238
rect 2672 1233 2677 1238
rect 2795 1235 2800 1240
rect 2818 1235 2823 1240
rect 2594 1225 2599 1230
rect 2730 1225 2735 1230
rect 2942 1235 2947 1240
rect 2965 1235 2970 1240
rect 2876 1227 2881 1232
rect 3023 1227 3028 1232
rect 484 1189 489 1194
rect 1872 1124 1877 1129
rect 1895 1124 1900 1129
rect 2016 1124 2021 1129
rect 2039 1124 2044 1129
rect 2165 1126 2170 1131
rect 2188 1126 2193 1131
rect 2310 1127 2315 1132
rect 2333 1127 2338 1132
rect 1953 1116 1958 1121
rect 2097 1116 2102 1121
rect 2246 1118 2251 1123
rect 2391 1119 2396 1124
rect 1565 1054 1570 1059
rect 1588 1054 1593 1059
rect 403 1028 408 1033
rect 421 1028 426 1033
rect 209 1010 214 1015
rect 269 1010 274 1015
rect 320 989 325 994
rect 338 989 343 994
rect 751 1012 756 1017
rect 774 1012 779 1017
rect 693 1004 698 1009
rect 898 1012 903 1017
rect 921 1012 926 1017
rect 1644 1047 1649 1052
rect 840 1004 845 1009
rect 1044 1010 1049 1015
rect 1067 1010 1072 1015
rect 986 1002 991 1007
rect 1180 1010 1185 1015
rect 1203 1010 1208 1015
rect 1122 1002 1127 1007
rect 481 967 486 972
rect 2273 944 2278 949
rect 2296 944 2301 949
rect 742 905 747 910
rect 765 905 770 910
rect 1564 936 1569 941
rect 1587 936 1592 941
rect 684 897 689 902
rect 887 904 892 909
rect 910 904 915 909
rect 1416 908 1421 913
rect 1454 908 1459 913
rect 1643 928 1648 933
rect 829 896 834 901
rect 1036 902 1041 907
rect 1059 902 1064 907
rect 978 894 983 899
rect 1180 902 1185 907
rect 1203 902 1208 907
rect 1122 894 1127 899
rect 2409 944 2414 949
rect 2432 944 2437 949
rect 2555 946 2560 951
rect 2578 946 2583 951
rect 2354 936 2359 941
rect 2490 936 2495 941
rect 2702 946 2707 951
rect 2725 946 2730 951
rect 2636 938 2641 943
rect 2783 938 2788 943
rect 18 837 23 842
rect 2081 875 2086 880
rect 406 843 411 848
rect 424 843 429 848
rect 2012 858 2017 863
rect 2036 858 2041 863
rect 1563 832 1568 837
rect 1586 832 1591 837
rect 2273 836 2278 841
rect 2296 836 2301 841
rect 77 821 82 826
rect 93 821 98 826
rect 109 821 114 826
rect 125 821 130 826
rect 212 825 217 830
rect 272 825 277 830
rect 323 804 328 809
rect 341 804 346 809
rect 1644 824 1649 829
rect 2417 836 2422 841
rect 2440 836 2445 841
rect 2566 838 2571 843
rect 2589 838 2594 843
rect 2711 839 2716 844
rect 2734 839 2739 844
rect 2354 828 2359 833
rect 2498 828 2503 833
rect 2647 830 2652 835
rect 2792 831 2797 836
rect 484 782 489 787
rect 1563 736 1568 741
rect 1586 736 1591 741
rect 1643 728 1648 733
rect 406 668 411 673
rect 424 668 429 673
rect 212 650 217 655
rect 272 650 277 655
rect 323 629 328 634
rect 341 629 346 634
rect 2162 638 2167 643
rect 2180 638 2185 643
rect 2024 620 2029 625
rect 484 607 489 612
rect 2079 599 2084 604
rect 2097 599 2102 604
rect 2240 577 2245 582
rect 1476 514 1481 519
rect 1539 496 1544 501
rect 1555 496 1560 501
rect 1571 496 1576 501
rect 2156 455 2161 460
rect 2174 455 2179 460
rect 2018 437 2023 442
rect 1360 389 1365 394
rect 1383 389 1388 394
rect 2073 416 2078 421
rect 2091 416 2096 421
rect 1302 381 1307 386
rect 1506 387 1511 392
rect 1529 387 1534 392
rect 1448 379 1453 384
rect 1642 387 1647 392
rect 1665 387 1670 392
rect 1584 379 1589 384
rect 2234 394 2239 399
rect 1310 266 1315 271
rect 1328 266 1333 271
rect 2144 283 2149 288
rect 2162 283 2167 288
rect 1648 266 1653 271
rect 1666 266 1671 271
rect 2006 265 2011 270
rect 1474 248 1479 253
rect 1393 227 1398 232
rect 1411 227 1416 232
rect 1806 248 1811 253
rect 2061 244 2066 249
rect 2079 244 2084 249
rect 1250 205 1255 210
rect 1588 205 1593 210
rect 1731 227 1736 232
rect 1749 227 1754 232
rect 2222 222 2227 227
rect 2135 99 2140 104
rect 2153 99 2158 104
rect 1997 81 2002 86
rect 2052 60 2057 65
rect 2070 60 2075 65
rect 2213 38 2218 43
rect 1444 -7 1449 -2
rect 1507 -25 1512 -20
rect 1523 -25 1528 -20
rect 1539 -25 1544 -20
rect 1328 -132 1333 -127
rect 1351 -132 1356 -127
rect 1270 -140 1275 -135
rect 1474 -134 1479 -129
rect 1497 -134 1502 -129
rect 1416 -142 1421 -137
rect 1610 -134 1615 -129
rect 1633 -134 1638 -129
rect 1552 -142 1557 -137
rect 1278 -255 1283 -250
rect 1296 -255 1301 -250
rect 1616 -255 1621 -250
rect 1634 -255 1639 -250
rect 1442 -273 1447 -268
rect 1218 -316 1223 -311
rect 1361 -294 1366 -289
rect 1379 -294 1384 -289
rect 1774 -273 1779 -268
rect 1556 -316 1561 -311
rect 1699 -294 1704 -289
rect 1717 -294 1722 -289
rect 1444 -458 1449 -453
rect 1507 -476 1512 -471
rect 1523 -476 1528 -471
rect 1539 -476 1544 -471
rect 1328 -583 1333 -578
rect 1351 -583 1356 -578
rect 1270 -591 1275 -586
rect 1474 -585 1479 -580
rect 1497 -585 1502 -580
rect 1416 -593 1421 -588
rect 1610 -585 1615 -580
rect 1633 -585 1638 -580
rect 1552 -593 1557 -588
rect 1278 -706 1283 -701
rect 1296 -706 1301 -701
rect 1616 -706 1621 -701
rect 1634 -706 1639 -701
rect 1442 -724 1447 -719
rect 1218 -767 1223 -762
rect 1361 -745 1366 -740
rect 1379 -745 1384 -740
rect 1774 -724 1779 -719
rect 1699 -745 1704 -740
rect 1717 -745 1722 -740
rect 1556 -767 1561 -762
rect 1435 -908 1440 -903
rect 1498 -926 1503 -921
rect 1514 -926 1519 -921
rect 1530 -926 1535 -921
rect 1319 -1033 1324 -1028
rect 1342 -1033 1347 -1028
rect 1261 -1041 1266 -1036
rect 1465 -1035 1470 -1030
rect 1488 -1035 1493 -1030
rect 1407 -1043 1412 -1038
rect 1601 -1035 1606 -1030
rect 1624 -1035 1629 -1030
rect 1543 -1043 1548 -1038
rect 1269 -1156 1274 -1151
rect 1287 -1156 1292 -1151
rect 1607 -1156 1612 -1151
rect 1625 -1156 1630 -1151
rect 1433 -1174 1438 -1169
rect 1352 -1195 1357 -1190
rect 1370 -1195 1375 -1190
rect 1765 -1174 1770 -1169
rect 1209 -1217 1214 -1212
rect 1547 -1217 1552 -1212
rect 1690 -1195 1695 -1190
rect 1708 -1195 1713 -1190
<< ptransistor >>
rect 936 1590 941 1595
rect 959 1590 964 1595
rect 878 1575 883 1580
rect 669 1489 674 1494
rect 685 1489 690 1494
rect 701 1489 706 1494
rect 717 1489 722 1494
rect 778 1493 783 1498
rect 835 1494 840 1499
rect 635 1290 640 1295
rect 690 1286 695 1291
rect 706 1286 711 1291
rect 722 1286 727 1291
rect 738 1286 743 1291
rect 754 1286 759 1291
rect 824 1290 829 1295
rect 212 1254 217 1259
rect 272 1254 277 1259
rect 883 1286 888 1291
rect 899 1286 904 1291
rect 915 1286 920 1291
rect 931 1286 936 1291
rect 982 1290 987 1295
rect 1045 1285 1050 1290
rect 1061 1285 1066 1290
rect 1077 1285 1082 1290
rect 1198 1287 1203 1292
rect 1221 1287 1226 1292
rect 323 1250 328 1255
rect 341 1250 346 1255
rect 1140 1272 1145 1277
rect 1872 1261 1877 1266
rect 1895 1261 1900 1266
rect 2008 1261 2013 1266
rect 2031 1261 2036 1266
rect 2154 1263 2159 1268
rect 2177 1263 2182 1268
rect 2301 1263 2306 1268
rect 2324 1263 2329 1268
rect 1953 1246 1958 1251
rect 2089 1246 2094 1251
rect 2235 1248 2240 1253
rect 2513 1262 2518 1267
rect 2536 1262 2541 1267
rect 2649 1262 2654 1267
rect 2672 1262 2677 1267
rect 2795 1264 2800 1269
rect 2818 1264 2823 1269
rect 2942 1264 2947 1269
rect 2965 1264 2970 1269
rect 2382 1248 2387 1253
rect 406 1211 411 1216
rect 424 1211 429 1216
rect 484 1211 489 1216
rect 2594 1247 2599 1252
rect 2730 1247 2735 1252
rect 2876 1249 2881 1254
rect 3023 1249 3028 1254
rect 1872 1153 1877 1158
rect 1895 1153 1900 1158
rect 2016 1153 2021 1158
rect 2039 1153 2044 1158
rect 2165 1155 2170 1160
rect 2188 1155 2193 1160
rect 2310 1156 2315 1161
rect 2333 1156 2338 1161
rect 1953 1138 1958 1143
rect 2097 1138 2102 1143
rect 2246 1140 2251 1145
rect 2391 1141 2396 1146
rect 1565 1083 1570 1088
rect 1588 1083 1593 1088
rect 209 1032 214 1037
rect 269 1032 274 1037
rect 1644 1069 1649 1074
rect 751 1041 756 1046
rect 774 1041 779 1046
rect 898 1041 903 1046
rect 921 1041 926 1046
rect 320 1028 325 1033
rect 338 1028 343 1033
rect 693 1026 698 1031
rect 840 1026 845 1031
rect 1044 1039 1049 1044
rect 1067 1039 1072 1044
rect 1180 1039 1185 1044
rect 1203 1039 1208 1044
rect 986 1024 991 1029
rect 403 989 408 994
rect 421 989 426 994
rect 481 989 486 994
rect 1122 1024 1127 1029
rect 2273 973 2278 978
rect 2296 973 2301 978
rect 2409 973 2414 978
rect 2432 973 2437 978
rect 2555 975 2560 980
rect 2578 975 2583 980
rect 2702 975 2707 980
rect 2725 975 2730 980
rect 1564 965 1569 970
rect 1587 965 1592 970
rect 742 934 747 939
rect 765 934 770 939
rect 684 919 689 924
rect 887 933 892 938
rect 910 933 915 938
rect 1643 950 1648 955
rect 2354 958 2359 963
rect 2490 958 2495 963
rect 2636 960 2641 965
rect 2783 960 2788 965
rect 829 918 834 923
rect 1036 931 1041 936
rect 1059 931 1064 936
rect 1180 931 1185 936
rect 1203 931 1208 936
rect 978 916 983 921
rect 1122 916 1127 921
rect 1416 930 1421 935
rect 1454 930 1459 935
rect 18 859 23 864
rect 2012 895 2017 900
rect 2036 895 2041 900
rect 2081 897 2086 902
rect 77 855 82 860
rect 93 855 98 860
rect 109 855 114 860
rect 125 855 130 860
rect 212 847 217 852
rect 272 847 277 852
rect 1563 861 1568 866
rect 1586 861 1591 866
rect 2273 865 2278 870
rect 2296 865 2301 870
rect 2417 865 2422 870
rect 2440 865 2445 870
rect 2566 867 2571 872
rect 2589 867 2594 872
rect 2711 868 2716 873
rect 2734 868 2739 873
rect 323 843 328 848
rect 341 843 346 848
rect 1644 846 1649 851
rect 2354 850 2359 855
rect 2498 850 2503 855
rect 2647 852 2652 857
rect 2792 853 2797 858
rect 406 804 411 809
rect 424 804 429 809
rect 484 804 489 809
rect 1563 765 1568 770
rect 1586 765 1591 770
rect 1643 750 1648 755
rect 212 672 217 677
rect 272 672 277 677
rect 323 668 328 673
rect 341 668 346 673
rect 2024 642 2029 647
rect 406 629 411 634
rect 424 629 429 634
rect 484 629 489 634
rect 2079 638 2084 643
rect 2097 638 2102 643
rect 2162 599 2167 604
rect 2180 599 2185 604
rect 2240 599 2245 604
rect 1476 536 1481 541
rect 1539 532 1544 537
rect 1555 532 1560 537
rect 1571 532 1576 537
rect 2018 459 2023 464
rect 2073 455 2078 460
rect 2091 455 2096 460
rect 1360 418 1365 423
rect 1383 418 1388 423
rect 1302 403 1307 408
rect 1506 416 1511 421
rect 1529 416 1534 421
rect 1642 416 1647 421
rect 1665 416 1670 421
rect 1448 401 1453 406
rect 1584 401 1589 406
rect 2156 416 2161 421
rect 2174 416 2179 421
rect 2234 416 2239 421
rect 1393 266 1398 271
rect 1411 266 1416 271
rect 1474 270 1479 275
rect 2006 287 2011 292
rect 2061 283 2066 288
rect 2079 283 2084 288
rect 1731 266 1736 271
rect 1749 266 1754 271
rect 1806 270 1811 275
rect 1250 227 1255 232
rect 1310 227 1315 232
rect 1328 227 1333 232
rect 1588 227 1593 232
rect 1648 227 1653 232
rect 1666 227 1671 232
rect 2144 244 2149 249
rect 2162 244 2167 249
rect 2222 244 2227 249
rect 1997 103 2002 108
rect 2052 99 2057 104
rect 2070 99 2075 104
rect 2135 60 2140 65
rect 2153 60 2158 65
rect 2213 60 2218 65
rect 1444 15 1449 20
rect 1507 11 1512 16
rect 1523 11 1528 16
rect 1539 11 1544 16
rect 1328 -103 1333 -98
rect 1351 -103 1356 -98
rect 1270 -118 1275 -113
rect 1474 -105 1479 -100
rect 1497 -105 1502 -100
rect 1610 -105 1615 -100
rect 1633 -105 1638 -100
rect 1416 -120 1421 -115
rect 1552 -120 1557 -115
rect 1361 -255 1366 -250
rect 1379 -255 1384 -250
rect 1442 -251 1447 -246
rect 1699 -255 1704 -250
rect 1717 -255 1722 -250
rect 1774 -251 1779 -246
rect 1218 -294 1223 -289
rect 1278 -294 1283 -289
rect 1296 -294 1301 -289
rect 1556 -294 1561 -289
rect 1616 -294 1621 -289
rect 1634 -294 1639 -289
rect 1444 -436 1449 -431
rect 1507 -440 1512 -435
rect 1523 -440 1528 -435
rect 1539 -440 1544 -435
rect 1328 -554 1333 -549
rect 1351 -554 1356 -549
rect 1270 -569 1275 -564
rect 1474 -556 1479 -551
rect 1497 -556 1502 -551
rect 1610 -556 1615 -551
rect 1633 -556 1638 -551
rect 1416 -571 1421 -566
rect 1552 -571 1557 -566
rect 1361 -706 1366 -701
rect 1379 -706 1384 -701
rect 1442 -702 1447 -697
rect 1699 -706 1704 -701
rect 1717 -706 1722 -701
rect 1774 -702 1779 -697
rect 1218 -745 1223 -740
rect 1278 -745 1283 -740
rect 1296 -745 1301 -740
rect 1556 -745 1561 -740
rect 1616 -745 1621 -740
rect 1634 -745 1639 -740
rect 1435 -886 1440 -881
rect 1498 -890 1503 -885
rect 1514 -890 1519 -885
rect 1530 -890 1535 -885
rect 1319 -1004 1324 -999
rect 1342 -1004 1347 -999
rect 1261 -1019 1266 -1014
rect 1465 -1006 1470 -1001
rect 1488 -1006 1493 -1001
rect 1601 -1006 1606 -1001
rect 1624 -1006 1629 -1001
rect 1407 -1021 1412 -1016
rect 1543 -1021 1548 -1016
rect 1352 -1156 1357 -1151
rect 1370 -1156 1375 -1151
rect 1433 -1152 1438 -1147
rect 1690 -1156 1695 -1151
rect 1708 -1156 1713 -1151
rect 1765 -1152 1770 -1147
rect 1209 -1195 1214 -1190
rect 1269 -1195 1274 -1190
rect 1287 -1195 1292 -1190
rect 1547 -1195 1552 -1190
rect 1607 -1195 1612 -1190
rect 1625 -1195 1630 -1190
<< ndiffusion >>
rect 934 1561 936 1566
rect 941 1561 943 1566
rect 957 1561 959 1566
rect 964 1561 966 1566
rect 875 1553 878 1558
rect 883 1553 885 1558
rect 776 1471 778 1476
rect 783 1471 786 1476
rect 833 1472 835 1477
rect 840 1472 843 1477
rect 666 1453 669 1458
rect 674 1453 677 1458
rect 682 1453 685 1458
rect 690 1453 693 1458
rect 698 1453 701 1458
rect 706 1453 709 1458
rect 714 1453 717 1458
rect 722 1453 725 1458
rect 632 1268 635 1273
rect 640 1268 642 1273
rect 821 1268 824 1273
rect 829 1268 831 1273
rect 979 1268 982 1273
rect 987 1268 989 1273
rect 403 1250 406 1255
rect 411 1250 424 1255
rect 429 1250 432 1255
rect 687 1252 690 1257
rect 695 1252 706 1257
rect 711 1252 722 1257
rect 727 1252 738 1257
rect 743 1252 754 1257
rect 759 1252 762 1257
rect 881 1252 883 1257
rect 888 1252 899 1257
rect 904 1252 915 1257
rect 920 1252 931 1257
rect 936 1252 939 1257
rect 210 1232 212 1237
rect 217 1232 220 1237
rect 269 1232 272 1237
rect 277 1232 279 1237
rect 1039 1251 1045 1256
rect 1050 1251 1061 1256
rect 1066 1251 1077 1256
rect 1082 1251 1085 1256
rect 1196 1258 1198 1263
rect 1203 1258 1205 1263
rect 1219 1258 1221 1263
rect 1226 1258 1228 1263
rect 1137 1250 1140 1255
rect 1145 1250 1147 1255
rect 1870 1232 1872 1237
rect 1877 1232 1879 1237
rect 1893 1232 1895 1237
rect 1900 1232 1902 1237
rect 320 1211 323 1216
rect 328 1211 341 1216
rect 346 1211 349 1216
rect 2006 1232 2008 1237
rect 2013 1232 2015 1237
rect 2029 1232 2031 1237
rect 2036 1232 2038 1237
rect 2152 1234 2154 1239
rect 2159 1234 2161 1239
rect 2175 1234 2177 1239
rect 2182 1234 2184 1239
rect 1951 1224 1953 1229
rect 1958 1224 1961 1229
rect 2087 1224 2089 1229
rect 2094 1224 2097 1229
rect 2299 1234 2301 1239
rect 2306 1234 2308 1239
rect 2322 1234 2324 1239
rect 2329 1234 2331 1239
rect 2233 1226 2235 1231
rect 2240 1226 2243 1231
rect 2511 1233 2513 1238
rect 2518 1233 2520 1238
rect 2534 1233 2536 1238
rect 2541 1233 2543 1238
rect 2380 1226 2382 1231
rect 2387 1226 2390 1231
rect 2647 1233 2649 1238
rect 2654 1233 2656 1238
rect 2670 1233 2672 1238
rect 2677 1233 2679 1238
rect 2793 1235 2795 1240
rect 2800 1235 2802 1240
rect 2816 1235 2818 1240
rect 2823 1235 2825 1240
rect 2592 1225 2594 1230
rect 2599 1225 2602 1230
rect 2728 1225 2730 1230
rect 2735 1225 2738 1230
rect 2940 1235 2942 1240
rect 2947 1235 2949 1240
rect 2963 1235 2965 1240
rect 2970 1235 2972 1240
rect 2874 1227 2876 1232
rect 2881 1227 2884 1232
rect 3021 1227 3023 1232
rect 3028 1227 3031 1232
rect 482 1189 484 1194
rect 489 1189 492 1194
rect 1870 1124 1872 1129
rect 1877 1124 1879 1129
rect 1893 1124 1895 1129
rect 1900 1124 1902 1129
rect 2014 1124 2016 1129
rect 2021 1124 2023 1129
rect 2037 1124 2039 1129
rect 2044 1124 2046 1129
rect 2163 1126 2165 1131
rect 2170 1126 2172 1131
rect 2186 1126 2188 1131
rect 2193 1126 2195 1131
rect 2308 1127 2310 1132
rect 2315 1127 2317 1132
rect 2331 1127 2333 1132
rect 2338 1127 2340 1132
rect 1951 1116 1953 1121
rect 1958 1116 1961 1121
rect 2095 1116 2097 1121
rect 2102 1116 2105 1121
rect 2244 1118 2246 1123
rect 2251 1118 2254 1123
rect 2389 1119 2391 1124
rect 2396 1119 2399 1124
rect 1563 1054 1565 1059
rect 1570 1054 1572 1059
rect 1586 1054 1588 1059
rect 1593 1054 1595 1059
rect 400 1028 403 1033
rect 408 1028 421 1033
rect 426 1028 429 1033
rect 207 1010 209 1015
rect 214 1010 217 1015
rect 266 1010 269 1015
rect 274 1010 276 1015
rect 317 989 320 994
rect 325 989 338 994
rect 343 989 346 994
rect 749 1012 751 1017
rect 756 1012 758 1017
rect 772 1012 774 1017
rect 779 1012 781 1017
rect 690 1004 693 1009
rect 698 1004 700 1009
rect 896 1012 898 1017
rect 903 1012 905 1017
rect 919 1012 921 1017
rect 926 1012 928 1017
rect 1642 1047 1644 1052
rect 1649 1047 1652 1052
rect 837 1004 840 1009
rect 845 1004 847 1009
rect 1042 1010 1044 1015
rect 1049 1010 1051 1015
rect 1065 1010 1067 1015
rect 1072 1010 1074 1015
rect 983 1002 986 1007
rect 991 1002 993 1007
rect 1178 1010 1180 1015
rect 1185 1010 1187 1015
rect 1201 1010 1203 1015
rect 1208 1010 1210 1015
rect 1119 1002 1122 1007
rect 1127 1002 1129 1007
rect 479 967 481 972
rect 486 967 489 972
rect 2271 944 2273 949
rect 2278 944 2280 949
rect 2294 944 2296 949
rect 2301 944 2303 949
rect 740 905 742 910
rect 747 905 749 910
rect 763 905 765 910
rect 770 905 772 910
rect 1562 936 1564 941
rect 1569 936 1571 941
rect 1585 936 1587 941
rect 1592 936 1594 941
rect 681 897 684 902
rect 689 897 691 902
rect 885 904 887 909
rect 892 904 894 909
rect 908 904 910 909
rect 915 904 917 909
rect 1414 908 1416 913
rect 1421 908 1424 913
rect 1452 908 1454 913
rect 1459 908 1462 913
rect 1641 928 1643 933
rect 1648 928 1651 933
rect 826 896 829 901
rect 834 896 836 901
rect 1034 902 1036 907
rect 1041 902 1043 907
rect 1057 902 1059 907
rect 1064 902 1066 907
rect 975 894 978 899
rect 983 894 985 899
rect 1178 902 1180 907
rect 1185 902 1187 907
rect 1201 902 1203 907
rect 1208 902 1210 907
rect 1119 894 1122 899
rect 1127 894 1129 899
rect 2407 944 2409 949
rect 2414 944 2416 949
rect 2430 944 2432 949
rect 2437 944 2439 949
rect 2553 946 2555 951
rect 2560 946 2562 951
rect 2576 946 2578 951
rect 2583 946 2585 951
rect 2352 936 2354 941
rect 2359 936 2362 941
rect 2488 936 2490 941
rect 2495 936 2498 941
rect 2700 946 2702 951
rect 2707 946 2709 951
rect 2723 946 2725 951
rect 2730 946 2732 951
rect 2634 938 2636 943
rect 2641 938 2644 943
rect 2781 938 2783 943
rect 2788 938 2791 943
rect 15 837 18 842
rect 23 837 25 842
rect 2079 875 2081 880
rect 2086 875 2089 880
rect 403 843 406 848
rect 411 843 424 848
rect 429 843 432 848
rect 2010 858 2012 863
rect 2017 858 2023 863
rect 2028 858 2036 863
rect 2041 858 2043 863
rect 1561 832 1563 837
rect 1568 832 1570 837
rect 1584 832 1586 837
rect 1591 832 1593 837
rect 2271 836 2273 841
rect 2278 836 2280 841
rect 2294 836 2296 841
rect 2301 836 2303 841
rect 75 821 77 826
rect 82 821 93 826
rect 98 821 109 826
rect 114 821 125 826
rect 130 821 133 826
rect 210 825 212 830
rect 217 825 220 830
rect 269 825 272 830
rect 277 825 279 830
rect 320 804 323 809
rect 328 804 341 809
rect 346 804 349 809
rect 1642 824 1644 829
rect 1649 824 1652 829
rect 2415 836 2417 841
rect 2422 836 2424 841
rect 2438 836 2440 841
rect 2445 836 2447 841
rect 2564 838 2566 843
rect 2571 838 2573 843
rect 2587 838 2589 843
rect 2594 838 2596 843
rect 2709 839 2711 844
rect 2716 839 2718 844
rect 2732 839 2734 844
rect 2739 839 2741 844
rect 2352 828 2354 833
rect 2359 828 2362 833
rect 2496 828 2498 833
rect 2503 828 2506 833
rect 2645 830 2647 835
rect 2652 830 2655 835
rect 2790 831 2792 836
rect 2797 831 2800 836
rect 482 782 484 787
rect 489 782 492 787
rect 1561 736 1563 741
rect 1568 736 1570 741
rect 1584 736 1586 741
rect 1591 736 1593 741
rect 1641 728 1643 733
rect 1648 728 1651 733
rect 403 668 406 673
rect 411 668 424 673
rect 429 668 432 673
rect 210 650 212 655
rect 217 650 220 655
rect 269 650 272 655
rect 277 650 279 655
rect 320 629 323 634
rect 328 629 341 634
rect 346 629 349 634
rect 2159 638 2162 643
rect 2167 638 2180 643
rect 2185 638 2188 643
rect 2021 620 2024 625
rect 2029 620 2031 625
rect 482 607 484 612
rect 489 607 492 612
rect 2076 599 2079 604
rect 2084 599 2097 604
rect 2102 599 2105 604
rect 2238 577 2240 582
rect 2245 577 2248 582
rect 1473 514 1476 519
rect 1481 514 1483 519
rect 1536 496 1539 501
rect 1544 496 1547 501
rect 1552 496 1555 501
rect 1560 496 1563 501
rect 1568 496 1571 501
rect 1576 496 1579 501
rect 2153 455 2156 460
rect 2161 455 2174 460
rect 2179 455 2182 460
rect 2015 437 2018 442
rect 2023 437 2025 442
rect 1358 389 1360 394
rect 1365 389 1367 394
rect 1381 389 1383 394
rect 1388 389 1390 394
rect 2070 416 2073 421
rect 2078 416 2091 421
rect 2096 416 2099 421
rect 1299 381 1302 386
rect 1307 381 1309 386
rect 1504 387 1506 392
rect 1511 387 1513 392
rect 1527 387 1529 392
rect 1534 387 1536 392
rect 1445 379 1448 384
rect 1453 379 1455 384
rect 1640 387 1642 392
rect 1647 387 1649 392
rect 1663 387 1665 392
rect 1670 387 1672 392
rect 1581 379 1584 384
rect 1589 379 1591 384
rect 2232 394 2234 399
rect 2239 394 2242 399
rect 1307 266 1310 271
rect 1315 266 1328 271
rect 1333 266 1336 271
rect 2141 283 2144 288
rect 2149 283 2162 288
rect 2167 283 2170 288
rect 1645 266 1648 271
rect 1653 266 1666 271
rect 1671 266 1674 271
rect 2003 265 2006 270
rect 2011 265 2013 270
rect 1472 248 1474 253
rect 1479 248 1482 253
rect 1390 227 1393 232
rect 1398 227 1411 232
rect 1416 227 1419 232
rect 1804 248 1806 253
rect 1811 248 1814 253
rect 2058 244 2061 249
rect 2066 244 2079 249
rect 2084 244 2087 249
rect 1247 205 1250 210
rect 1255 205 1257 210
rect 1585 205 1588 210
rect 1593 205 1595 210
rect 1728 227 1731 232
rect 1736 227 1749 232
rect 1754 227 1757 232
rect 2220 222 2222 227
rect 2227 222 2230 227
rect 2132 99 2135 104
rect 2140 99 2153 104
rect 2158 99 2161 104
rect 1994 81 1997 86
rect 2002 81 2004 86
rect 2049 60 2052 65
rect 2057 60 2070 65
rect 2075 60 2078 65
rect 2211 38 2213 43
rect 2218 38 2221 43
rect 1441 -7 1444 -2
rect 1449 -7 1451 -2
rect 1504 -25 1507 -20
rect 1512 -25 1515 -20
rect 1520 -25 1523 -20
rect 1528 -25 1531 -20
rect 1536 -25 1539 -20
rect 1544 -25 1547 -20
rect 1326 -132 1328 -127
rect 1333 -132 1335 -127
rect 1349 -132 1351 -127
rect 1356 -132 1358 -127
rect 1267 -140 1270 -135
rect 1275 -140 1277 -135
rect 1472 -134 1474 -129
rect 1479 -134 1481 -129
rect 1495 -134 1497 -129
rect 1502 -134 1504 -129
rect 1413 -142 1416 -137
rect 1421 -142 1423 -137
rect 1608 -134 1610 -129
rect 1615 -134 1617 -129
rect 1631 -134 1633 -129
rect 1638 -134 1640 -129
rect 1549 -142 1552 -137
rect 1557 -142 1559 -137
rect 1275 -255 1278 -250
rect 1283 -255 1296 -250
rect 1301 -255 1304 -250
rect 1613 -255 1616 -250
rect 1621 -255 1634 -250
rect 1639 -255 1642 -250
rect 1440 -273 1442 -268
rect 1447 -273 1450 -268
rect 1215 -316 1218 -311
rect 1223 -316 1225 -311
rect 1358 -294 1361 -289
rect 1366 -294 1379 -289
rect 1384 -294 1387 -289
rect 1772 -273 1774 -268
rect 1779 -273 1782 -268
rect 1553 -316 1556 -311
rect 1561 -316 1563 -311
rect 1696 -294 1699 -289
rect 1704 -294 1717 -289
rect 1722 -294 1725 -289
rect 1441 -458 1444 -453
rect 1449 -458 1451 -453
rect 1504 -476 1507 -471
rect 1512 -476 1515 -471
rect 1520 -476 1523 -471
rect 1528 -476 1531 -471
rect 1536 -476 1539 -471
rect 1544 -476 1547 -471
rect 1326 -583 1328 -578
rect 1333 -583 1335 -578
rect 1349 -583 1351 -578
rect 1356 -583 1358 -578
rect 1267 -591 1270 -586
rect 1275 -591 1277 -586
rect 1472 -585 1474 -580
rect 1479 -585 1481 -580
rect 1495 -585 1497 -580
rect 1502 -585 1504 -580
rect 1413 -593 1416 -588
rect 1421 -593 1423 -588
rect 1608 -585 1610 -580
rect 1615 -585 1617 -580
rect 1631 -585 1633 -580
rect 1638 -585 1640 -580
rect 1549 -593 1552 -588
rect 1557 -593 1559 -588
rect 1275 -706 1278 -701
rect 1283 -706 1296 -701
rect 1301 -706 1304 -701
rect 1613 -706 1616 -701
rect 1621 -706 1634 -701
rect 1639 -706 1642 -701
rect 1440 -724 1442 -719
rect 1447 -724 1450 -719
rect 1215 -767 1218 -762
rect 1223 -767 1225 -762
rect 1358 -745 1361 -740
rect 1366 -745 1379 -740
rect 1384 -745 1387 -740
rect 1772 -724 1774 -719
rect 1779 -724 1782 -719
rect 1696 -745 1699 -740
rect 1704 -745 1717 -740
rect 1722 -745 1725 -740
rect 1553 -767 1556 -762
rect 1561 -767 1563 -762
rect 1432 -908 1435 -903
rect 1440 -908 1442 -903
rect 1495 -926 1498 -921
rect 1503 -926 1506 -921
rect 1511 -926 1514 -921
rect 1519 -926 1522 -921
rect 1527 -926 1530 -921
rect 1535 -926 1538 -921
rect 1317 -1033 1319 -1028
rect 1324 -1033 1326 -1028
rect 1340 -1033 1342 -1028
rect 1347 -1033 1349 -1028
rect 1258 -1041 1261 -1036
rect 1266 -1041 1268 -1036
rect 1463 -1035 1465 -1030
rect 1470 -1035 1472 -1030
rect 1486 -1035 1488 -1030
rect 1493 -1035 1495 -1030
rect 1404 -1043 1407 -1038
rect 1412 -1043 1414 -1038
rect 1599 -1035 1601 -1030
rect 1606 -1035 1608 -1030
rect 1622 -1035 1624 -1030
rect 1629 -1035 1631 -1030
rect 1540 -1043 1543 -1038
rect 1548 -1043 1550 -1038
rect 1266 -1156 1269 -1151
rect 1274 -1156 1287 -1151
rect 1292 -1156 1295 -1151
rect 1604 -1156 1607 -1151
rect 1612 -1156 1625 -1151
rect 1630 -1156 1633 -1151
rect 1431 -1174 1433 -1169
rect 1438 -1174 1441 -1169
rect 1349 -1195 1352 -1190
rect 1357 -1195 1370 -1190
rect 1375 -1195 1378 -1190
rect 1763 -1174 1765 -1169
rect 1770 -1174 1773 -1169
rect 1206 -1217 1209 -1212
rect 1214 -1217 1216 -1212
rect 1544 -1217 1547 -1212
rect 1552 -1217 1554 -1212
rect 1687 -1195 1690 -1190
rect 1695 -1195 1708 -1190
rect 1713 -1195 1716 -1190
<< pdiffusion >>
rect 934 1590 936 1595
rect 941 1590 947 1595
rect 952 1590 959 1595
rect 964 1590 966 1595
rect 875 1575 878 1580
rect 883 1575 885 1580
rect 666 1489 669 1494
rect 674 1489 685 1494
rect 690 1489 701 1494
rect 706 1489 717 1494
rect 722 1489 725 1494
rect 776 1493 778 1498
rect 783 1493 786 1498
rect 833 1494 835 1499
rect 840 1494 843 1499
rect 632 1290 635 1295
rect 640 1290 642 1295
rect 687 1286 690 1291
rect 695 1286 698 1291
rect 703 1286 706 1291
rect 711 1286 714 1291
rect 719 1286 722 1291
rect 727 1286 730 1291
rect 735 1286 738 1291
rect 743 1286 746 1291
rect 751 1286 754 1291
rect 759 1286 762 1291
rect 821 1290 824 1295
rect 829 1290 831 1295
rect 210 1254 212 1259
rect 217 1254 220 1259
rect 269 1254 272 1259
rect 277 1254 279 1259
rect 880 1286 883 1291
rect 888 1286 891 1291
rect 896 1286 899 1291
rect 904 1286 907 1291
rect 912 1286 915 1291
rect 920 1286 923 1291
rect 928 1286 931 1291
rect 936 1286 939 1291
rect 979 1290 982 1295
rect 987 1290 989 1295
rect 1042 1285 1045 1290
rect 1050 1285 1053 1290
rect 1058 1285 1061 1290
rect 1066 1285 1069 1290
rect 1074 1285 1077 1290
rect 1082 1285 1085 1290
rect 1196 1287 1198 1292
rect 1203 1287 1209 1292
rect 1214 1287 1221 1292
rect 1226 1287 1228 1292
rect 320 1250 323 1255
rect 328 1250 341 1255
rect 346 1250 349 1255
rect 1137 1272 1140 1277
rect 1145 1272 1147 1277
rect 1870 1261 1872 1266
rect 1877 1261 1884 1266
rect 1889 1261 1895 1266
rect 1900 1261 1902 1266
rect 2006 1261 2008 1266
rect 2013 1261 2020 1266
rect 2025 1261 2031 1266
rect 2036 1261 2038 1266
rect 2152 1263 2154 1268
rect 2159 1263 2166 1268
rect 2171 1263 2177 1268
rect 2182 1263 2184 1268
rect 2299 1263 2301 1268
rect 2306 1263 2313 1268
rect 2318 1263 2324 1268
rect 2329 1263 2331 1268
rect 1951 1246 1953 1251
rect 1958 1246 1961 1251
rect 2087 1246 2089 1251
rect 2094 1246 2097 1251
rect 2233 1248 2235 1253
rect 2240 1248 2243 1253
rect 2511 1262 2513 1267
rect 2518 1262 2525 1267
rect 2530 1262 2536 1267
rect 2541 1262 2543 1267
rect 2647 1262 2649 1267
rect 2654 1262 2661 1267
rect 2666 1262 2672 1267
rect 2677 1262 2679 1267
rect 2793 1264 2795 1269
rect 2800 1264 2807 1269
rect 2812 1264 2818 1269
rect 2823 1264 2825 1269
rect 2940 1264 2942 1269
rect 2947 1264 2954 1269
rect 2959 1264 2965 1269
rect 2970 1264 2972 1269
rect 2380 1248 2382 1253
rect 2387 1248 2390 1253
rect 403 1211 406 1216
rect 411 1211 424 1216
rect 429 1211 432 1216
rect 482 1211 484 1216
rect 489 1211 492 1216
rect 2592 1247 2594 1252
rect 2599 1247 2602 1252
rect 2728 1247 2730 1252
rect 2735 1247 2738 1252
rect 2874 1249 2876 1254
rect 2881 1249 2884 1254
rect 3021 1249 3023 1254
rect 3028 1249 3031 1254
rect 1870 1153 1872 1158
rect 1877 1153 1884 1158
rect 1889 1153 1895 1158
rect 1900 1153 1902 1158
rect 2014 1153 2016 1158
rect 2021 1153 2028 1158
rect 2033 1153 2039 1158
rect 2044 1153 2046 1158
rect 2163 1155 2165 1160
rect 2170 1155 2177 1160
rect 2182 1155 2188 1160
rect 2193 1155 2195 1160
rect 2308 1156 2310 1161
rect 2315 1156 2322 1161
rect 2327 1156 2333 1161
rect 2338 1156 2340 1161
rect 1951 1138 1953 1143
rect 1958 1138 1961 1143
rect 2095 1138 2097 1143
rect 2102 1138 2105 1143
rect 2244 1140 2246 1145
rect 2251 1140 2254 1145
rect 2389 1141 2391 1146
rect 2396 1141 2399 1146
rect 1563 1083 1565 1088
rect 1570 1083 1577 1088
rect 1582 1083 1588 1088
rect 1593 1083 1595 1088
rect 207 1032 209 1037
rect 214 1032 217 1037
rect 266 1032 269 1037
rect 274 1032 276 1037
rect 1642 1069 1644 1074
rect 1649 1069 1652 1074
rect 749 1041 751 1046
rect 756 1041 762 1046
rect 767 1041 774 1046
rect 779 1041 781 1046
rect 896 1041 898 1046
rect 903 1041 909 1046
rect 914 1041 921 1046
rect 926 1041 928 1046
rect 317 1028 320 1033
rect 325 1028 338 1033
rect 343 1028 346 1033
rect 690 1026 693 1031
rect 698 1026 700 1031
rect 837 1026 840 1031
rect 845 1026 847 1031
rect 1042 1039 1044 1044
rect 1049 1039 1055 1044
rect 1060 1039 1067 1044
rect 1072 1039 1074 1044
rect 1178 1039 1180 1044
rect 1185 1039 1191 1044
rect 1196 1039 1203 1044
rect 1208 1039 1210 1044
rect 983 1024 986 1029
rect 991 1024 993 1029
rect 400 989 403 994
rect 408 989 421 994
rect 426 989 429 994
rect 479 989 481 994
rect 486 989 489 994
rect 1119 1024 1122 1029
rect 1127 1024 1129 1029
rect 2271 973 2273 978
rect 2278 973 2285 978
rect 2290 973 2296 978
rect 2301 973 2303 978
rect 2407 973 2409 978
rect 2414 973 2421 978
rect 2426 973 2432 978
rect 2437 973 2439 978
rect 2553 975 2555 980
rect 2560 975 2567 980
rect 2572 975 2578 980
rect 2583 975 2585 980
rect 2700 975 2702 980
rect 2707 975 2714 980
rect 2719 975 2725 980
rect 2730 975 2732 980
rect 1562 965 1564 970
rect 1569 965 1576 970
rect 1581 965 1587 970
rect 1592 965 1594 970
rect 740 934 742 939
rect 747 934 753 939
rect 758 934 765 939
rect 770 934 772 939
rect 681 919 684 924
rect 689 919 691 924
rect 885 933 887 938
rect 892 933 898 938
rect 903 933 910 938
rect 915 933 917 938
rect 1641 950 1643 955
rect 1648 950 1651 955
rect 2352 958 2354 963
rect 2359 958 2362 963
rect 2488 958 2490 963
rect 2495 958 2498 963
rect 2634 960 2636 965
rect 2641 960 2644 965
rect 2781 960 2783 965
rect 2788 960 2791 965
rect 826 918 829 923
rect 834 918 836 923
rect 1034 931 1036 936
rect 1041 931 1047 936
rect 1052 931 1059 936
rect 1064 931 1066 936
rect 1178 931 1180 936
rect 1185 931 1191 936
rect 1196 931 1203 936
rect 1208 931 1210 936
rect 975 916 978 921
rect 983 916 985 921
rect 1119 916 1122 921
rect 1127 916 1129 921
rect 1414 930 1416 935
rect 1421 930 1424 935
rect 1452 930 1454 935
rect 1459 930 1462 935
rect 15 859 18 864
rect 23 859 25 864
rect 2010 895 2012 900
rect 2017 895 2019 900
rect 2034 895 2036 900
rect 2041 895 2043 900
rect 2079 897 2081 902
rect 2086 897 2089 902
rect 74 855 77 860
rect 82 855 85 860
rect 90 855 93 860
rect 98 855 101 860
rect 106 855 109 860
rect 114 855 117 860
rect 122 855 125 860
rect 130 855 133 860
rect 210 847 212 852
rect 217 847 220 852
rect 269 847 272 852
rect 277 847 279 852
rect 1561 861 1563 866
rect 1568 861 1575 866
rect 1580 861 1586 866
rect 1591 861 1593 866
rect 2271 865 2273 870
rect 2278 865 2285 870
rect 2290 865 2296 870
rect 2301 865 2303 870
rect 2415 865 2417 870
rect 2422 865 2429 870
rect 2434 865 2440 870
rect 2445 865 2447 870
rect 2564 867 2566 872
rect 2571 867 2578 872
rect 2583 867 2589 872
rect 2594 867 2596 872
rect 2709 868 2711 873
rect 2716 868 2723 873
rect 2728 868 2734 873
rect 2739 868 2741 873
rect 320 843 323 848
rect 328 843 341 848
rect 346 843 349 848
rect 1642 846 1644 851
rect 1649 846 1652 851
rect 2352 850 2354 855
rect 2359 850 2362 855
rect 2496 850 2498 855
rect 2503 850 2506 855
rect 2645 852 2647 857
rect 2652 852 2655 857
rect 2790 853 2792 858
rect 2797 853 2800 858
rect 403 804 406 809
rect 411 804 424 809
rect 429 804 432 809
rect 482 804 484 809
rect 489 804 492 809
rect 1561 765 1563 770
rect 1568 765 1575 770
rect 1580 765 1586 770
rect 1591 765 1593 770
rect 1641 750 1643 755
rect 1648 750 1651 755
rect 210 672 212 677
rect 217 672 220 677
rect 269 672 272 677
rect 277 672 279 677
rect 320 668 323 673
rect 328 668 341 673
rect 346 668 349 673
rect 2021 642 2024 647
rect 2029 642 2031 647
rect 403 629 406 634
rect 411 629 424 634
rect 429 629 432 634
rect 482 629 484 634
rect 489 629 492 634
rect 2076 638 2079 643
rect 2084 638 2097 643
rect 2102 638 2105 643
rect 2159 599 2162 604
rect 2167 599 2180 604
rect 2185 599 2188 604
rect 2238 599 2240 604
rect 2245 599 2248 604
rect 1473 536 1476 541
rect 1481 536 1483 541
rect 1536 532 1539 537
rect 1544 532 1555 537
rect 1560 532 1571 537
rect 1576 532 1579 537
rect 2015 459 2018 464
rect 2023 459 2025 464
rect 2070 455 2073 460
rect 2078 455 2091 460
rect 2096 455 2099 460
rect 1358 418 1360 423
rect 1365 418 1371 423
rect 1376 418 1383 423
rect 1388 418 1390 423
rect 1299 403 1302 408
rect 1307 403 1309 408
rect 1504 416 1506 421
rect 1511 416 1517 421
rect 1522 416 1529 421
rect 1534 416 1536 421
rect 1640 416 1642 421
rect 1647 416 1653 421
rect 1658 416 1665 421
rect 1670 416 1672 421
rect 1445 401 1448 406
rect 1453 401 1455 406
rect 1581 401 1584 406
rect 1589 401 1591 406
rect 2153 416 2156 421
rect 2161 416 2174 421
rect 2179 416 2182 421
rect 2232 416 2234 421
rect 2239 416 2242 421
rect 1390 266 1393 271
rect 1398 266 1411 271
rect 1416 266 1419 271
rect 1472 270 1474 275
rect 1479 270 1482 275
rect 2003 287 2006 292
rect 2011 287 2013 292
rect 2058 283 2061 288
rect 2066 283 2079 288
rect 2084 283 2087 288
rect 1728 266 1731 271
rect 1736 266 1749 271
rect 1754 266 1757 271
rect 1804 270 1806 275
rect 1811 270 1814 275
rect 1247 227 1250 232
rect 1255 227 1257 232
rect 1307 227 1310 232
rect 1315 227 1328 232
rect 1333 227 1336 232
rect 1585 227 1588 232
rect 1593 227 1595 232
rect 1645 227 1648 232
rect 1653 227 1666 232
rect 1671 227 1674 232
rect 2141 244 2144 249
rect 2149 244 2162 249
rect 2167 244 2170 249
rect 2220 244 2222 249
rect 2227 244 2230 249
rect 1994 103 1997 108
rect 2002 103 2004 108
rect 2049 99 2052 104
rect 2057 99 2070 104
rect 2075 99 2078 104
rect 2132 60 2135 65
rect 2140 60 2153 65
rect 2158 60 2161 65
rect 2211 60 2213 65
rect 2218 60 2221 65
rect 1441 15 1444 20
rect 1449 15 1451 20
rect 1504 11 1507 16
rect 1512 11 1523 16
rect 1528 11 1539 16
rect 1544 11 1547 16
rect 1326 -103 1328 -98
rect 1333 -103 1339 -98
rect 1344 -103 1351 -98
rect 1356 -103 1358 -98
rect 1267 -118 1270 -113
rect 1275 -118 1277 -113
rect 1472 -105 1474 -100
rect 1479 -105 1485 -100
rect 1490 -105 1497 -100
rect 1502 -105 1504 -100
rect 1608 -105 1610 -100
rect 1615 -105 1621 -100
rect 1626 -105 1633 -100
rect 1638 -105 1640 -100
rect 1413 -120 1416 -115
rect 1421 -120 1423 -115
rect 1549 -120 1552 -115
rect 1557 -120 1559 -115
rect 1358 -255 1361 -250
rect 1366 -255 1379 -250
rect 1384 -255 1387 -250
rect 1440 -251 1442 -246
rect 1447 -251 1450 -246
rect 1696 -255 1699 -250
rect 1704 -255 1717 -250
rect 1722 -255 1725 -250
rect 1772 -251 1774 -246
rect 1779 -251 1782 -246
rect 1215 -294 1218 -289
rect 1223 -294 1225 -289
rect 1275 -294 1278 -289
rect 1283 -294 1296 -289
rect 1301 -294 1304 -289
rect 1553 -294 1556 -289
rect 1561 -294 1563 -289
rect 1613 -294 1616 -289
rect 1621 -294 1634 -289
rect 1639 -294 1642 -289
rect 1441 -436 1444 -431
rect 1449 -436 1451 -431
rect 1504 -440 1507 -435
rect 1512 -440 1523 -435
rect 1528 -440 1539 -435
rect 1544 -440 1547 -435
rect 1326 -554 1328 -549
rect 1333 -554 1339 -549
rect 1344 -554 1351 -549
rect 1356 -554 1358 -549
rect 1267 -569 1270 -564
rect 1275 -569 1277 -564
rect 1472 -556 1474 -551
rect 1479 -556 1485 -551
rect 1490 -556 1497 -551
rect 1502 -556 1504 -551
rect 1608 -556 1610 -551
rect 1615 -556 1621 -551
rect 1626 -556 1633 -551
rect 1638 -556 1640 -551
rect 1413 -571 1416 -566
rect 1421 -571 1423 -566
rect 1549 -571 1552 -566
rect 1557 -571 1559 -566
rect 1358 -706 1361 -701
rect 1366 -706 1379 -701
rect 1384 -706 1387 -701
rect 1440 -702 1442 -697
rect 1447 -702 1450 -697
rect 1696 -706 1699 -701
rect 1704 -706 1717 -701
rect 1722 -706 1725 -701
rect 1772 -702 1774 -697
rect 1779 -702 1782 -697
rect 1215 -745 1218 -740
rect 1223 -745 1225 -740
rect 1275 -745 1278 -740
rect 1283 -745 1296 -740
rect 1301 -745 1304 -740
rect 1553 -745 1556 -740
rect 1561 -745 1563 -740
rect 1613 -745 1616 -740
rect 1621 -745 1634 -740
rect 1639 -745 1642 -740
rect 1432 -886 1435 -881
rect 1440 -886 1442 -881
rect 1495 -890 1498 -885
rect 1503 -890 1514 -885
rect 1519 -890 1530 -885
rect 1535 -890 1538 -885
rect 1317 -1004 1319 -999
rect 1324 -1004 1330 -999
rect 1335 -1004 1342 -999
rect 1347 -1004 1349 -999
rect 1258 -1019 1261 -1014
rect 1266 -1019 1268 -1014
rect 1463 -1006 1465 -1001
rect 1470 -1006 1476 -1001
rect 1481 -1006 1488 -1001
rect 1493 -1006 1495 -1001
rect 1599 -1006 1601 -1001
rect 1606 -1006 1612 -1001
rect 1617 -1006 1624 -1001
rect 1629 -1006 1631 -1001
rect 1404 -1021 1407 -1016
rect 1412 -1021 1414 -1016
rect 1540 -1021 1543 -1016
rect 1548 -1021 1550 -1016
rect 1349 -1156 1352 -1151
rect 1357 -1156 1370 -1151
rect 1375 -1156 1378 -1151
rect 1431 -1152 1433 -1147
rect 1438 -1152 1441 -1147
rect 1687 -1156 1690 -1151
rect 1695 -1156 1708 -1151
rect 1713 -1156 1716 -1151
rect 1763 -1152 1765 -1147
rect 1770 -1152 1773 -1147
rect 1206 -1195 1209 -1190
rect 1214 -1195 1216 -1190
rect 1266 -1195 1269 -1190
rect 1274 -1195 1287 -1190
rect 1292 -1195 1295 -1190
rect 1544 -1195 1547 -1190
rect 1552 -1195 1554 -1190
rect 1604 -1195 1607 -1190
rect 1612 -1195 1625 -1190
rect 1630 -1195 1633 -1190
<< ndcontact >>
rect 929 1561 934 1566
rect 943 1561 947 1566
rect 953 1561 957 1566
rect 966 1561 971 1566
rect 870 1553 875 1558
rect 885 1553 890 1558
rect 771 1471 776 1476
rect 786 1471 791 1476
rect 828 1472 833 1477
rect 843 1472 848 1477
rect 661 1453 666 1458
rect 677 1453 682 1458
rect 693 1453 698 1458
rect 709 1453 714 1458
rect 725 1453 730 1458
rect 627 1268 632 1273
rect 642 1268 647 1273
rect 816 1268 821 1273
rect 831 1268 836 1273
rect 974 1268 979 1273
rect 989 1268 994 1273
rect 398 1250 403 1255
rect 432 1250 437 1255
rect 682 1252 687 1257
rect 762 1252 767 1257
rect 876 1252 881 1257
rect 939 1252 944 1257
rect 205 1232 210 1237
rect 220 1232 225 1237
rect 264 1232 269 1237
rect 279 1232 284 1237
rect 1034 1251 1039 1256
rect 1085 1251 1090 1256
rect 1191 1258 1196 1263
rect 1205 1258 1209 1263
rect 1215 1258 1219 1263
rect 1228 1258 1233 1263
rect 1132 1250 1137 1255
rect 1147 1250 1152 1255
rect 1865 1232 1870 1237
rect 1879 1232 1883 1237
rect 1889 1232 1893 1237
rect 1902 1232 1907 1237
rect 315 1211 320 1216
rect 349 1211 354 1216
rect 2001 1232 2006 1237
rect 2015 1232 2019 1237
rect 2025 1232 2029 1237
rect 2038 1232 2043 1237
rect 2147 1234 2152 1239
rect 2161 1234 2165 1239
rect 2171 1234 2175 1239
rect 2184 1234 2189 1239
rect 1946 1224 1951 1229
rect 1961 1224 1966 1229
rect 2082 1224 2087 1229
rect 2097 1224 2102 1229
rect 2294 1234 2299 1239
rect 2308 1234 2312 1239
rect 2318 1234 2322 1239
rect 2331 1234 2336 1239
rect 2228 1226 2233 1231
rect 2243 1226 2248 1231
rect 2506 1233 2511 1238
rect 2520 1233 2524 1238
rect 2530 1233 2534 1238
rect 2543 1233 2548 1238
rect 2375 1226 2380 1231
rect 2390 1226 2395 1231
rect 2642 1233 2647 1238
rect 2656 1233 2660 1238
rect 2666 1233 2670 1238
rect 2679 1233 2684 1238
rect 2788 1235 2793 1240
rect 2802 1235 2806 1240
rect 2812 1235 2816 1240
rect 2825 1235 2830 1240
rect 2587 1225 2592 1230
rect 2602 1225 2607 1230
rect 2723 1225 2728 1230
rect 2738 1225 2743 1230
rect 2935 1235 2940 1240
rect 2949 1235 2953 1240
rect 2959 1235 2963 1240
rect 2972 1235 2977 1240
rect 2869 1227 2874 1232
rect 2884 1227 2889 1232
rect 3016 1227 3021 1232
rect 3031 1227 3036 1232
rect 477 1189 482 1194
rect 492 1189 497 1194
rect 1865 1124 1870 1129
rect 1879 1124 1883 1129
rect 1889 1124 1893 1129
rect 1902 1124 1907 1129
rect 2009 1124 2014 1129
rect 2023 1124 2027 1129
rect 2033 1124 2037 1129
rect 2046 1124 2051 1129
rect 2158 1126 2163 1131
rect 2172 1126 2176 1131
rect 2182 1126 2186 1131
rect 2195 1126 2200 1131
rect 2303 1127 2308 1132
rect 2317 1127 2321 1132
rect 2327 1127 2331 1132
rect 2340 1127 2345 1132
rect 1946 1116 1951 1121
rect 1961 1116 1966 1121
rect 2090 1116 2095 1121
rect 2105 1116 2110 1121
rect 2239 1118 2244 1123
rect 2254 1118 2259 1123
rect 2384 1119 2389 1124
rect 2399 1119 2404 1124
rect 1558 1054 1563 1059
rect 1572 1054 1576 1059
rect 1582 1054 1586 1059
rect 1595 1054 1600 1059
rect 395 1028 400 1033
rect 429 1028 434 1033
rect 202 1010 207 1015
rect 217 1010 222 1015
rect 261 1010 266 1015
rect 276 1010 281 1015
rect 312 989 317 994
rect 346 989 351 994
rect 744 1012 749 1017
rect 758 1012 762 1017
rect 768 1012 772 1017
rect 781 1012 786 1017
rect 685 1004 690 1009
rect 700 1004 705 1009
rect 891 1012 896 1017
rect 905 1012 909 1017
rect 915 1012 919 1017
rect 928 1012 933 1017
rect 1637 1047 1642 1052
rect 1652 1047 1657 1052
rect 832 1004 837 1009
rect 847 1004 852 1009
rect 1037 1010 1042 1015
rect 1051 1010 1055 1015
rect 1061 1010 1065 1015
rect 1074 1010 1079 1015
rect 978 1002 983 1007
rect 993 1002 998 1007
rect 1173 1010 1178 1015
rect 1187 1010 1191 1015
rect 1197 1010 1201 1015
rect 1210 1010 1215 1015
rect 1114 1002 1119 1007
rect 1129 1002 1134 1007
rect 474 967 479 972
rect 489 967 494 972
rect 2266 944 2271 949
rect 2280 944 2284 949
rect 2290 944 2294 949
rect 2303 944 2308 949
rect 735 905 740 910
rect 749 905 753 910
rect 759 905 763 910
rect 772 905 777 910
rect 1557 936 1562 941
rect 1571 936 1575 941
rect 1581 936 1585 941
rect 1594 936 1599 941
rect 676 897 681 902
rect 691 897 696 902
rect 880 904 885 909
rect 894 904 898 909
rect 904 904 908 909
rect 917 904 922 909
rect 1409 908 1414 913
rect 1424 908 1429 913
rect 1447 908 1452 913
rect 1462 908 1467 913
rect 1636 928 1641 933
rect 1651 928 1656 933
rect 821 896 826 901
rect 836 896 841 901
rect 1029 902 1034 907
rect 1043 902 1047 907
rect 1053 902 1057 907
rect 1066 902 1071 907
rect 970 894 975 899
rect 985 894 990 899
rect 1173 902 1178 907
rect 1187 902 1191 907
rect 1197 902 1201 907
rect 1210 902 1215 907
rect 1114 894 1119 899
rect 1129 894 1134 899
rect 2402 944 2407 949
rect 2416 944 2420 949
rect 2426 944 2430 949
rect 2439 944 2444 949
rect 2548 946 2553 951
rect 2562 946 2566 951
rect 2572 946 2576 951
rect 2585 946 2590 951
rect 2347 936 2352 941
rect 2362 936 2367 941
rect 2483 936 2488 941
rect 2498 936 2503 941
rect 2695 946 2700 951
rect 2709 946 2713 951
rect 2719 946 2723 951
rect 2732 946 2737 951
rect 2629 938 2634 943
rect 2644 938 2649 943
rect 2776 938 2781 943
rect 2791 938 2796 943
rect 10 837 15 842
rect 25 837 30 842
rect 2074 875 2079 880
rect 2089 875 2094 880
rect 398 843 403 848
rect 432 843 437 848
rect 2005 858 2010 863
rect 2023 858 2028 863
rect 2043 858 2048 863
rect 1556 832 1561 837
rect 1570 832 1574 837
rect 1580 832 1584 837
rect 1593 832 1598 837
rect 2266 836 2271 841
rect 2280 836 2284 841
rect 2290 836 2294 841
rect 2303 836 2308 841
rect 70 821 75 826
rect 133 821 138 826
rect 205 825 210 830
rect 220 825 225 830
rect 264 825 269 830
rect 279 825 284 830
rect 315 804 320 809
rect 349 804 354 809
rect 1637 824 1642 829
rect 1652 824 1657 829
rect 2410 836 2415 841
rect 2424 836 2428 841
rect 2434 836 2438 841
rect 2447 836 2452 841
rect 2559 838 2564 843
rect 2573 838 2577 843
rect 2583 838 2587 843
rect 2596 838 2601 843
rect 2704 839 2709 844
rect 2718 839 2722 844
rect 2728 839 2732 844
rect 2741 839 2746 844
rect 2347 828 2352 833
rect 2362 828 2367 833
rect 2491 828 2496 833
rect 2506 828 2511 833
rect 2640 830 2645 835
rect 2655 830 2660 835
rect 2785 831 2790 836
rect 2800 831 2805 836
rect 477 782 482 787
rect 492 782 497 787
rect 1556 736 1561 741
rect 1570 736 1574 741
rect 1580 736 1584 741
rect 1593 736 1598 741
rect 1636 728 1641 733
rect 1651 728 1656 733
rect 398 668 403 673
rect 432 668 437 673
rect 205 650 210 655
rect 220 650 225 655
rect 264 650 269 655
rect 279 650 284 655
rect 315 629 320 634
rect 349 629 354 634
rect 2154 638 2159 643
rect 2188 638 2193 643
rect 2016 620 2021 625
rect 2031 620 2036 625
rect 477 607 482 612
rect 492 607 497 612
rect 2071 599 2076 604
rect 2105 599 2110 604
rect 2233 577 2238 582
rect 2248 577 2253 582
rect 1468 514 1473 519
rect 1483 514 1488 519
rect 1531 496 1536 501
rect 1547 496 1552 501
rect 1563 496 1568 501
rect 1579 496 1584 501
rect 2148 455 2153 460
rect 2182 455 2187 460
rect 2010 437 2015 442
rect 2025 437 2030 442
rect 1353 389 1358 394
rect 1367 389 1371 394
rect 1377 389 1381 394
rect 1390 389 1395 394
rect 2065 416 2070 421
rect 2099 416 2104 421
rect 1294 381 1299 386
rect 1309 381 1314 386
rect 1499 387 1504 392
rect 1513 387 1517 392
rect 1523 387 1527 392
rect 1536 387 1541 392
rect 1440 379 1445 384
rect 1455 379 1460 384
rect 1635 387 1640 392
rect 1649 387 1653 392
rect 1659 387 1663 392
rect 1672 387 1677 392
rect 1576 379 1581 384
rect 1591 379 1596 384
rect 2227 394 2232 399
rect 2242 394 2247 399
rect 1302 266 1307 271
rect 1336 266 1341 271
rect 2136 283 2141 288
rect 2170 283 2175 288
rect 1640 266 1645 271
rect 1674 266 1679 271
rect 1998 265 2003 270
rect 2013 265 2018 270
rect 1467 248 1472 253
rect 1482 248 1487 253
rect 1385 227 1390 232
rect 1419 227 1424 232
rect 1799 248 1804 253
rect 1814 248 1819 253
rect 2053 244 2058 249
rect 2087 244 2092 249
rect 1242 205 1247 210
rect 1257 205 1262 210
rect 1580 205 1585 210
rect 1595 205 1600 210
rect 1723 227 1728 232
rect 1757 227 1762 232
rect 2215 222 2220 227
rect 2230 222 2235 227
rect 2127 99 2132 104
rect 2161 99 2166 104
rect 1989 81 1994 86
rect 2004 81 2009 86
rect 2044 60 2049 65
rect 2078 60 2083 65
rect 2206 38 2211 43
rect 2221 38 2226 43
rect 1436 -7 1441 -2
rect 1451 -7 1456 -2
rect 1499 -25 1504 -20
rect 1515 -25 1520 -20
rect 1531 -25 1536 -20
rect 1547 -25 1552 -20
rect 1321 -132 1326 -127
rect 1335 -132 1339 -127
rect 1345 -132 1349 -127
rect 1358 -132 1363 -127
rect 1262 -140 1267 -135
rect 1277 -140 1282 -135
rect 1467 -134 1472 -129
rect 1481 -134 1485 -129
rect 1491 -134 1495 -129
rect 1504 -134 1509 -129
rect 1408 -142 1413 -137
rect 1423 -142 1428 -137
rect 1603 -134 1608 -129
rect 1617 -134 1621 -129
rect 1627 -134 1631 -129
rect 1640 -134 1645 -129
rect 1544 -142 1549 -137
rect 1559 -142 1564 -137
rect 1270 -255 1275 -250
rect 1304 -255 1309 -250
rect 1608 -255 1613 -250
rect 1642 -255 1647 -250
rect 1435 -273 1440 -268
rect 1450 -273 1455 -268
rect 1210 -316 1215 -311
rect 1225 -316 1230 -311
rect 1353 -294 1358 -289
rect 1387 -294 1392 -289
rect 1767 -273 1772 -268
rect 1782 -273 1787 -268
rect 1548 -316 1553 -311
rect 1563 -316 1568 -311
rect 1691 -294 1696 -289
rect 1725 -294 1730 -289
rect 1436 -458 1441 -453
rect 1451 -458 1456 -453
rect 1499 -476 1504 -471
rect 1515 -476 1520 -471
rect 1531 -476 1536 -471
rect 1547 -476 1552 -471
rect 1321 -583 1326 -578
rect 1335 -583 1339 -578
rect 1345 -583 1349 -578
rect 1358 -583 1363 -578
rect 1262 -591 1267 -586
rect 1277 -591 1282 -586
rect 1467 -585 1472 -580
rect 1481 -585 1485 -580
rect 1491 -585 1495 -580
rect 1504 -585 1509 -580
rect 1408 -593 1413 -588
rect 1423 -593 1428 -588
rect 1603 -585 1608 -580
rect 1617 -585 1621 -580
rect 1627 -585 1631 -580
rect 1640 -585 1645 -580
rect 1544 -593 1549 -588
rect 1559 -593 1564 -588
rect 1270 -706 1275 -701
rect 1304 -706 1309 -701
rect 1608 -706 1613 -701
rect 1642 -706 1647 -701
rect 1435 -724 1440 -719
rect 1450 -724 1455 -719
rect 1210 -767 1215 -762
rect 1225 -767 1230 -762
rect 1353 -745 1358 -740
rect 1387 -745 1392 -740
rect 1767 -724 1772 -719
rect 1782 -724 1787 -719
rect 1691 -745 1696 -740
rect 1725 -745 1730 -740
rect 1548 -767 1553 -762
rect 1563 -767 1568 -762
rect 1427 -908 1432 -903
rect 1442 -908 1447 -903
rect 1490 -926 1495 -921
rect 1506 -926 1511 -921
rect 1522 -926 1527 -921
rect 1538 -926 1543 -921
rect 1312 -1033 1317 -1028
rect 1326 -1033 1330 -1028
rect 1336 -1033 1340 -1028
rect 1349 -1033 1354 -1028
rect 1253 -1041 1258 -1036
rect 1268 -1041 1273 -1036
rect 1458 -1035 1463 -1030
rect 1472 -1035 1476 -1030
rect 1482 -1035 1486 -1030
rect 1495 -1035 1500 -1030
rect 1399 -1043 1404 -1038
rect 1414 -1043 1419 -1038
rect 1594 -1035 1599 -1030
rect 1608 -1035 1612 -1030
rect 1618 -1035 1622 -1030
rect 1631 -1035 1636 -1030
rect 1535 -1043 1540 -1038
rect 1550 -1043 1555 -1038
rect 1261 -1156 1266 -1151
rect 1295 -1156 1300 -1151
rect 1599 -1156 1604 -1151
rect 1633 -1156 1638 -1151
rect 1426 -1174 1431 -1169
rect 1441 -1174 1446 -1169
rect 1344 -1195 1349 -1190
rect 1378 -1195 1383 -1190
rect 1758 -1174 1763 -1169
rect 1773 -1174 1778 -1169
rect 1201 -1217 1206 -1212
rect 1216 -1217 1221 -1212
rect 1539 -1217 1544 -1212
rect 1554 -1217 1559 -1212
rect 1682 -1195 1687 -1190
rect 1716 -1195 1721 -1190
<< pdcontact >>
rect 929 1590 934 1595
rect 947 1590 952 1595
rect 966 1590 971 1595
rect 870 1575 875 1580
rect 885 1575 890 1580
rect 661 1489 666 1494
rect 725 1489 730 1494
rect 771 1493 776 1498
rect 786 1493 791 1498
rect 828 1494 833 1499
rect 843 1494 848 1499
rect 627 1290 632 1295
rect 642 1290 647 1295
rect 682 1286 687 1291
rect 698 1286 703 1291
rect 714 1286 719 1291
rect 730 1286 735 1291
rect 746 1286 751 1291
rect 762 1286 767 1291
rect 816 1290 821 1295
rect 831 1290 836 1295
rect 205 1254 210 1259
rect 220 1254 225 1259
rect 264 1254 269 1259
rect 279 1254 284 1259
rect 875 1286 880 1291
rect 891 1286 896 1291
rect 907 1286 912 1291
rect 923 1286 928 1291
rect 939 1286 944 1291
rect 974 1290 979 1295
rect 989 1290 994 1295
rect 1037 1285 1042 1290
rect 1053 1285 1058 1290
rect 1069 1285 1074 1290
rect 1085 1285 1090 1290
rect 1191 1287 1196 1292
rect 1209 1287 1214 1292
rect 1228 1287 1233 1292
rect 315 1250 320 1255
rect 349 1250 354 1255
rect 1132 1272 1137 1277
rect 1147 1272 1152 1277
rect 1865 1261 1870 1266
rect 1884 1261 1889 1266
rect 1902 1261 1907 1266
rect 2001 1261 2006 1266
rect 2020 1261 2025 1266
rect 2038 1261 2043 1266
rect 2147 1263 2152 1268
rect 2166 1263 2171 1268
rect 2184 1263 2189 1268
rect 2294 1263 2299 1268
rect 2313 1263 2318 1268
rect 2331 1263 2336 1268
rect 1946 1246 1951 1251
rect 1961 1246 1966 1251
rect 2082 1246 2087 1251
rect 2097 1246 2102 1251
rect 2228 1248 2233 1253
rect 2243 1248 2248 1253
rect 2506 1262 2511 1267
rect 2525 1262 2530 1267
rect 2543 1262 2548 1267
rect 2642 1262 2647 1267
rect 2661 1262 2666 1267
rect 2679 1262 2684 1267
rect 2788 1264 2793 1269
rect 2807 1264 2812 1269
rect 2825 1264 2830 1269
rect 2935 1264 2940 1269
rect 2954 1264 2959 1269
rect 2972 1264 2977 1269
rect 2375 1248 2380 1253
rect 2390 1248 2395 1253
rect 398 1211 403 1216
rect 432 1211 437 1216
rect 477 1211 482 1216
rect 492 1211 497 1216
rect 2587 1247 2592 1252
rect 2602 1247 2607 1252
rect 2723 1247 2728 1252
rect 2738 1247 2743 1252
rect 2869 1249 2874 1254
rect 2884 1249 2889 1254
rect 3016 1249 3021 1254
rect 3031 1249 3036 1254
rect 1865 1153 1870 1158
rect 1884 1153 1889 1158
rect 1902 1153 1907 1158
rect 2009 1153 2014 1158
rect 2028 1153 2033 1158
rect 2046 1153 2051 1158
rect 2158 1155 2163 1160
rect 2177 1155 2182 1160
rect 2195 1155 2200 1160
rect 2303 1156 2308 1161
rect 2322 1156 2327 1161
rect 2340 1156 2345 1161
rect 1946 1138 1951 1143
rect 1961 1138 1966 1143
rect 2090 1138 2095 1143
rect 2105 1138 2110 1143
rect 2239 1140 2244 1145
rect 2254 1140 2259 1145
rect 2384 1141 2389 1146
rect 2399 1141 2404 1146
rect 1558 1083 1563 1088
rect 1577 1083 1582 1088
rect 1595 1083 1600 1088
rect 202 1032 207 1037
rect 217 1032 222 1037
rect 261 1032 266 1037
rect 276 1032 281 1037
rect 1637 1069 1642 1074
rect 1652 1069 1657 1074
rect 744 1041 749 1046
rect 762 1041 767 1046
rect 781 1041 786 1046
rect 891 1041 896 1046
rect 909 1041 914 1046
rect 928 1041 933 1046
rect 312 1028 317 1033
rect 346 1028 351 1033
rect 685 1026 690 1031
rect 700 1026 705 1031
rect 832 1026 837 1031
rect 847 1026 852 1031
rect 1037 1039 1042 1044
rect 1055 1039 1060 1044
rect 1074 1039 1079 1044
rect 1173 1039 1178 1044
rect 1191 1039 1196 1044
rect 1210 1039 1215 1044
rect 978 1024 983 1029
rect 993 1024 998 1029
rect 395 989 400 994
rect 429 989 434 994
rect 474 989 479 994
rect 489 989 494 994
rect 1114 1024 1119 1029
rect 1129 1024 1134 1029
rect 2266 973 2271 978
rect 2285 973 2290 978
rect 2303 973 2308 978
rect 2402 973 2407 978
rect 2421 973 2426 978
rect 2439 973 2444 978
rect 2548 975 2553 980
rect 2567 975 2572 980
rect 2585 975 2590 980
rect 2695 975 2700 980
rect 2714 975 2719 980
rect 2732 975 2737 980
rect 1557 965 1562 970
rect 1576 965 1581 970
rect 1594 965 1599 970
rect 735 934 740 939
rect 753 934 758 939
rect 772 934 777 939
rect 676 919 681 924
rect 691 919 696 924
rect 880 933 885 938
rect 898 933 903 938
rect 917 933 922 938
rect 1636 950 1641 955
rect 1651 950 1656 955
rect 2347 958 2352 963
rect 2362 958 2367 963
rect 2483 958 2488 963
rect 2498 958 2503 963
rect 2629 960 2634 965
rect 2644 960 2649 965
rect 2776 960 2781 965
rect 2791 960 2796 965
rect 821 918 826 923
rect 836 918 841 923
rect 1029 931 1034 936
rect 1047 931 1052 936
rect 1066 931 1071 936
rect 1173 931 1178 936
rect 1191 931 1196 936
rect 1210 931 1215 936
rect 970 916 975 921
rect 985 916 990 921
rect 1114 916 1119 921
rect 1129 916 1134 921
rect 1409 930 1414 935
rect 1424 930 1429 935
rect 1447 930 1452 935
rect 1462 930 1467 935
rect 10 859 15 864
rect 25 859 30 864
rect 2005 895 2010 900
rect 2019 895 2024 900
rect 2029 895 2034 900
rect 2043 895 2048 900
rect 2074 897 2079 902
rect 2089 897 2094 902
rect 69 855 74 860
rect 85 855 90 860
rect 101 855 106 860
rect 117 855 122 860
rect 133 855 138 860
rect 205 847 210 852
rect 220 847 225 852
rect 264 847 269 852
rect 279 847 284 852
rect 1556 861 1561 866
rect 1575 861 1580 866
rect 1593 861 1598 866
rect 2266 865 2271 870
rect 2285 865 2290 870
rect 2303 865 2308 870
rect 2410 865 2415 870
rect 2429 865 2434 870
rect 2447 865 2452 870
rect 2559 867 2564 872
rect 2578 867 2583 872
rect 2596 867 2601 872
rect 2704 868 2709 873
rect 2723 868 2728 873
rect 2741 868 2746 873
rect 315 843 320 848
rect 349 843 354 848
rect 1637 846 1642 851
rect 1652 846 1657 851
rect 2347 850 2352 855
rect 2362 850 2367 855
rect 2491 850 2496 855
rect 2506 850 2511 855
rect 2640 852 2645 857
rect 2655 852 2660 857
rect 2785 853 2790 858
rect 2800 853 2805 858
rect 398 804 403 809
rect 432 804 437 809
rect 477 804 482 809
rect 492 804 497 809
rect 1556 765 1561 770
rect 1575 765 1580 770
rect 1593 765 1598 770
rect 1636 750 1641 755
rect 1651 750 1656 755
rect 205 672 210 677
rect 220 672 225 677
rect 264 672 269 677
rect 279 672 284 677
rect 315 668 320 673
rect 349 668 354 673
rect 2016 642 2021 647
rect 2031 642 2036 647
rect 398 629 403 634
rect 432 629 437 634
rect 477 629 482 634
rect 492 629 497 634
rect 2071 638 2076 643
rect 2105 638 2110 643
rect 2154 599 2159 604
rect 2188 599 2193 604
rect 2233 599 2238 604
rect 2248 599 2253 604
rect 1468 536 1473 541
rect 1483 536 1488 541
rect 1531 532 1536 537
rect 1579 532 1584 537
rect 2010 459 2015 464
rect 2025 459 2030 464
rect 2065 455 2070 460
rect 2099 455 2104 460
rect 1353 418 1358 423
rect 1371 418 1376 423
rect 1390 418 1395 423
rect 1294 403 1299 408
rect 1309 403 1314 408
rect 1499 416 1504 421
rect 1517 416 1522 421
rect 1536 416 1541 421
rect 1635 416 1640 421
rect 1653 416 1658 421
rect 1672 416 1677 421
rect 1440 401 1445 406
rect 1455 401 1460 406
rect 1576 401 1581 406
rect 1591 401 1596 406
rect 2148 416 2153 421
rect 2182 416 2187 421
rect 2227 416 2232 421
rect 2242 416 2247 421
rect 1385 266 1390 271
rect 1419 266 1424 271
rect 1467 270 1472 275
rect 1482 270 1487 275
rect 1998 287 2003 292
rect 2013 287 2018 292
rect 2053 283 2058 288
rect 2087 283 2092 288
rect 1723 266 1728 271
rect 1757 266 1762 271
rect 1799 270 1804 275
rect 1814 270 1819 275
rect 1242 227 1247 232
rect 1257 227 1262 232
rect 1302 227 1307 232
rect 1336 227 1341 232
rect 1580 227 1585 232
rect 1595 227 1600 232
rect 1640 227 1645 232
rect 1674 227 1679 232
rect 2136 244 2141 249
rect 2170 244 2175 249
rect 2215 244 2220 249
rect 2230 244 2235 249
rect 1989 103 1994 108
rect 2004 103 2009 108
rect 2044 99 2049 104
rect 2078 99 2083 104
rect 2127 60 2132 65
rect 2161 60 2166 65
rect 2206 60 2211 65
rect 2221 60 2226 65
rect 1436 15 1441 20
rect 1451 15 1456 20
rect 1499 11 1504 16
rect 1547 11 1552 16
rect 1321 -103 1326 -98
rect 1339 -103 1344 -98
rect 1358 -103 1363 -98
rect 1262 -118 1267 -113
rect 1277 -118 1282 -113
rect 1467 -105 1472 -100
rect 1485 -105 1490 -100
rect 1504 -105 1509 -100
rect 1603 -105 1608 -100
rect 1621 -105 1626 -100
rect 1640 -105 1645 -100
rect 1408 -120 1413 -115
rect 1423 -120 1428 -115
rect 1544 -120 1549 -115
rect 1559 -120 1564 -115
rect 1353 -255 1358 -250
rect 1387 -255 1392 -250
rect 1435 -251 1440 -246
rect 1450 -251 1455 -246
rect 1691 -255 1696 -250
rect 1725 -255 1730 -250
rect 1767 -251 1772 -246
rect 1782 -251 1787 -246
rect 1210 -294 1215 -289
rect 1225 -294 1230 -289
rect 1270 -294 1275 -289
rect 1304 -294 1309 -289
rect 1548 -294 1553 -289
rect 1563 -294 1568 -289
rect 1608 -294 1613 -289
rect 1642 -294 1647 -289
rect 1436 -436 1441 -431
rect 1451 -436 1456 -431
rect 1499 -440 1504 -435
rect 1547 -440 1552 -435
rect 1321 -554 1326 -549
rect 1339 -554 1344 -549
rect 1358 -554 1363 -549
rect 1262 -569 1267 -564
rect 1277 -569 1282 -564
rect 1467 -556 1472 -551
rect 1485 -556 1490 -551
rect 1504 -556 1509 -551
rect 1603 -556 1608 -551
rect 1621 -556 1626 -551
rect 1640 -556 1645 -551
rect 1408 -571 1413 -566
rect 1423 -571 1428 -566
rect 1544 -571 1549 -566
rect 1559 -571 1564 -566
rect 1353 -706 1358 -701
rect 1387 -706 1392 -701
rect 1435 -702 1440 -697
rect 1450 -702 1455 -697
rect 1691 -706 1696 -701
rect 1725 -706 1730 -701
rect 1767 -702 1772 -697
rect 1782 -702 1787 -697
rect 1210 -745 1215 -740
rect 1225 -745 1230 -740
rect 1270 -745 1275 -740
rect 1304 -745 1309 -740
rect 1548 -745 1553 -740
rect 1563 -745 1568 -740
rect 1608 -745 1613 -740
rect 1642 -745 1647 -740
rect 1427 -886 1432 -881
rect 1442 -886 1447 -881
rect 1490 -890 1495 -885
rect 1538 -890 1543 -885
rect 1312 -1004 1317 -999
rect 1330 -1004 1335 -999
rect 1349 -1004 1354 -999
rect 1253 -1019 1258 -1014
rect 1268 -1019 1273 -1014
rect 1458 -1006 1463 -1001
rect 1476 -1006 1481 -1001
rect 1495 -1006 1500 -1001
rect 1594 -1006 1599 -1001
rect 1612 -1006 1617 -1001
rect 1631 -1006 1636 -1001
rect 1399 -1021 1404 -1016
rect 1414 -1021 1419 -1016
rect 1535 -1021 1540 -1016
rect 1550 -1021 1555 -1016
rect 1344 -1156 1349 -1151
rect 1378 -1156 1383 -1151
rect 1426 -1152 1431 -1147
rect 1441 -1152 1446 -1147
rect 1682 -1156 1687 -1151
rect 1716 -1156 1721 -1151
rect 1758 -1152 1763 -1147
rect 1773 -1152 1778 -1147
rect 1201 -1195 1206 -1190
rect 1216 -1195 1221 -1190
rect 1261 -1195 1266 -1190
rect 1295 -1195 1300 -1190
rect 1539 -1195 1544 -1190
rect 1554 -1195 1559 -1190
rect 1599 -1195 1604 -1190
rect 1633 -1195 1638 -1190
<< nsubstratencontact >>
rect 975 1590 980 1595
rect 897 1575 902 1580
rect 737 1489 742 1494
rect 759 1493 764 1498
rect 816 1494 821 1499
rect 654 1290 659 1295
rect 843 1290 848 1295
rect 193 1254 198 1259
rect 291 1254 296 1259
rect 863 1286 868 1291
rect 1001 1290 1006 1295
rect 1027 1285 1032 1290
rect 1237 1287 1242 1292
rect 303 1250 308 1255
rect 1159 1272 1164 1277
rect 1856 1261 1861 1266
rect 1992 1261 1997 1266
rect 2139 1263 2143 1268
rect 2285 1263 2290 1268
rect 1934 1246 1939 1251
rect 2070 1246 2075 1251
rect 2216 1248 2221 1253
rect 2497 1262 2502 1267
rect 2633 1262 2638 1267
rect 2779 1264 2784 1269
rect 2926 1264 2931 1269
rect 2363 1248 2368 1253
rect 383 1209 389 1215
rect 465 1211 470 1216
rect 2575 1247 2580 1252
rect 2711 1247 2716 1252
rect 2857 1249 2862 1254
rect 3004 1249 3009 1254
rect 1856 1153 1861 1158
rect 2000 1153 2005 1158
rect 2149 1155 2154 1160
rect 2294 1156 2299 1161
rect 1934 1138 1939 1143
rect 2078 1138 2083 1143
rect 2227 1140 2232 1145
rect 2372 1141 2377 1146
rect 1549 1083 1554 1088
rect 190 1032 195 1037
rect 288 1032 293 1037
rect 1625 1069 1630 1074
rect 790 1041 795 1046
rect 937 1041 942 1046
rect 300 1028 305 1033
rect 712 1026 717 1031
rect 859 1026 864 1031
rect 1083 1039 1088 1044
rect 1219 1039 1224 1044
rect 1005 1024 1010 1029
rect 380 990 386 995
rect 462 989 467 994
rect 1141 1024 1146 1029
rect 2257 973 2262 978
rect 2393 973 2398 978
rect 2539 975 2544 980
rect 2686 975 2691 980
rect 1548 965 1553 970
rect 781 934 786 939
rect 703 919 708 924
rect 926 933 931 938
rect 1624 950 1629 955
rect 2335 958 2340 963
rect 2471 958 2476 963
rect 2617 960 2622 965
rect 2764 960 2769 965
rect 848 918 853 923
rect 1075 931 1080 936
rect 1219 931 1224 936
rect 997 916 1002 921
rect 1141 916 1146 921
rect 1397 930 1402 935
rect 37 859 42 864
rect 1995 895 2000 900
rect 2062 897 2067 902
rect 57 855 62 860
rect 168 847 173 852
rect 291 847 296 852
rect 1547 861 1552 866
rect 2257 865 2262 870
rect 2401 865 2406 870
rect 2550 867 2555 872
rect 2695 868 2700 873
rect 303 843 308 848
rect 1625 846 1630 851
rect 2335 850 2340 855
rect 2479 850 2484 855
rect 2628 852 2633 857
rect 2773 853 2778 858
rect 383 802 388 808
rect 465 804 470 809
rect 1547 765 1552 770
rect 1624 750 1629 755
rect 193 672 198 677
rect 291 672 296 677
rect 303 668 308 673
rect 2043 642 2048 647
rect 383 629 388 634
rect 465 629 470 634
rect 2059 638 2064 643
rect 2139 597 2144 602
rect 2221 599 2226 604
rect 1495 536 1500 541
rect 1522 532 1527 537
rect 2053 455 2058 460
rect 1399 418 1404 423
rect 1321 403 1326 408
rect 1545 416 1550 421
rect 1681 416 1686 421
rect 1467 401 1472 406
rect 1603 401 1608 406
rect 2133 414 2139 420
rect 2215 416 2220 421
rect 1431 266 1436 271
rect 1455 270 1460 275
rect 2041 283 2046 288
rect 1769 266 1774 271
rect 1787 270 1792 275
rect 1269 227 1274 232
rect 1347 228 1354 235
rect 1607 227 1612 232
rect 1689 225 1694 231
rect 2121 242 2126 247
rect 2203 244 2208 249
rect 2032 99 2037 104
rect 2112 62 2117 67
rect 2194 60 2199 65
rect 1463 15 1468 20
rect 1490 11 1495 16
rect 1367 -103 1372 -98
rect 1289 -118 1294 -113
rect 1513 -105 1518 -100
rect 1649 -105 1654 -100
rect 1435 -120 1440 -115
rect 1571 -120 1576 -115
rect 1399 -255 1404 -250
rect 1423 -251 1428 -246
rect 1737 -255 1742 -250
rect 1755 -251 1760 -246
rect 1237 -294 1242 -289
rect 1319 -296 1324 -291
rect 1575 -294 1580 -289
rect 1657 -296 1663 -290
rect 1463 -436 1468 -431
rect 1490 -440 1495 -435
rect 1367 -554 1372 -549
rect 1289 -569 1294 -564
rect 1513 -556 1518 -551
rect 1649 -556 1654 -551
rect 1435 -571 1440 -566
rect 1571 -571 1576 -566
rect 1399 -706 1404 -701
rect 1423 -702 1428 -697
rect 1737 -706 1742 -701
rect 1755 -702 1760 -697
rect 1237 -745 1242 -740
rect 1319 -747 1324 -742
rect 1575 -745 1580 -740
rect 1655 -744 1661 -738
rect 1454 -886 1459 -881
rect 1481 -890 1486 -885
rect 1358 -1004 1363 -999
rect 1280 -1019 1285 -1014
rect 1504 -1006 1509 -1001
rect 1640 -1006 1645 -1001
rect 1426 -1021 1431 -1016
rect 1562 -1021 1567 -1016
rect 1390 -1156 1395 -1151
rect 1414 -1152 1419 -1147
rect 1728 -1156 1733 -1151
rect 1746 -1152 1751 -1147
rect 1228 -1195 1233 -1190
rect 1308 -1195 1312 -1190
rect 1566 -1195 1571 -1190
rect 1648 -1197 1654 -1192
<< polysilicon >>
rect 936 1595 941 1609
rect 959 1595 964 1609
rect 878 1580 883 1583
rect 878 1566 883 1575
rect 936 1566 941 1590
rect 959 1566 964 1590
rect 878 1562 882 1566
rect 878 1558 883 1562
rect 878 1548 883 1553
rect 936 1542 941 1561
rect 959 1542 964 1561
rect 778 1498 783 1501
rect 835 1499 840 1502
rect 669 1494 674 1497
rect 685 1494 690 1497
rect 701 1494 706 1497
rect 717 1494 722 1497
rect 669 1458 674 1489
rect 685 1458 690 1489
rect 701 1458 706 1489
rect 717 1458 722 1489
rect 778 1484 783 1493
rect 835 1485 840 1494
rect 779 1480 783 1484
rect 836 1481 840 1485
rect 778 1476 783 1480
rect 835 1477 840 1481
rect 778 1466 783 1471
rect 835 1467 840 1472
rect 669 1442 674 1453
rect 685 1442 690 1453
rect 701 1442 706 1453
rect 717 1443 722 1453
rect 635 1295 640 1298
rect 690 1291 695 1295
rect 706 1291 711 1295
rect 722 1291 727 1310
rect 738 1291 743 1310
rect 824 1295 829 1298
rect 754 1291 759 1295
rect 635 1281 640 1290
rect 883 1291 888 1310
rect 899 1291 904 1310
rect 915 1291 920 1295
rect 931 1291 936 1310
rect 982 1295 987 1298
rect 341 1276 379 1277
rect 635 1277 639 1281
rect 384 1276 429 1277
rect 341 1272 429 1276
rect 635 1273 640 1277
rect 212 1259 217 1262
rect 272 1259 277 1262
rect 323 1255 328 1259
rect 341 1255 346 1272
rect 406 1255 411 1259
rect 424 1255 429 1272
rect 635 1263 640 1268
rect 690 1257 695 1286
rect 706 1257 711 1286
rect 722 1257 727 1286
rect 738 1257 743 1286
rect 754 1257 759 1286
rect 824 1281 829 1290
rect 1045 1290 1050 1295
rect 1061 1290 1066 1312
rect 1077 1290 1082 1310
rect 1198 1292 1203 1306
rect 1221 1292 1226 1306
rect 824 1277 828 1281
rect 824 1273 829 1277
rect 824 1263 829 1268
rect 883 1257 888 1286
rect 899 1257 904 1286
rect 915 1257 920 1286
rect 931 1257 936 1286
rect 982 1281 987 1290
rect 982 1277 986 1281
rect 982 1273 987 1277
rect 982 1263 987 1268
rect 212 1245 217 1254
rect 213 1241 217 1245
rect 212 1237 217 1241
rect 272 1245 277 1254
rect 1045 1256 1050 1285
rect 1061 1256 1066 1285
rect 1077 1256 1082 1285
rect 1140 1277 1145 1280
rect 1140 1263 1145 1272
rect 1198 1263 1203 1287
rect 1221 1263 1226 1287
rect 1872 1266 1877 1280
rect 1895 1266 1900 1280
rect 2008 1266 2013 1280
rect 2031 1266 2036 1280
rect 2154 1268 2159 1282
rect 2177 1268 2182 1282
rect 2301 1268 2306 1282
rect 2324 1268 2329 1282
rect 1140 1259 1144 1263
rect 272 1241 276 1245
rect 272 1237 277 1241
rect 323 1238 328 1250
rect 341 1246 346 1250
rect 406 1238 411 1250
rect 424 1246 429 1250
rect 324 1233 346 1238
rect 406 1233 429 1238
rect 690 1233 695 1252
rect 212 1227 217 1232
rect 272 1227 277 1232
rect 304 1221 328 1226
rect 304 1213 309 1221
rect 323 1216 328 1221
rect 341 1216 346 1233
rect 406 1216 411 1220
rect 424 1216 429 1233
rect 706 1232 711 1252
rect 722 1235 727 1252
rect 738 1235 743 1252
rect 754 1232 759 1252
rect 883 1245 888 1252
rect 899 1245 904 1252
rect 915 1235 920 1252
rect 931 1235 936 1252
rect 1140 1255 1145 1259
rect 2513 1267 2518 1281
rect 2536 1267 2541 1281
rect 2649 1267 2654 1281
rect 2672 1267 2677 1281
rect 2795 1269 2800 1283
rect 2818 1269 2823 1283
rect 2942 1269 2947 1283
rect 2965 1269 2970 1283
rect 1045 1236 1050 1251
rect 1061 1237 1066 1251
rect 1077 1237 1082 1251
rect 1140 1245 1145 1250
rect 1198 1239 1203 1258
rect 1221 1239 1226 1258
rect 1872 1237 1877 1261
rect 1895 1237 1900 1261
rect 1953 1251 1958 1254
rect 1953 1237 1958 1246
rect 2008 1237 2013 1261
rect 2031 1237 2036 1261
rect 2089 1251 2094 1254
rect 2089 1237 2094 1246
rect 2154 1239 2159 1263
rect 2177 1239 2182 1263
rect 2235 1253 2240 1256
rect 2235 1239 2240 1248
rect 2301 1239 2306 1263
rect 2324 1239 2329 1263
rect 2382 1253 2387 1256
rect 2382 1239 2387 1248
rect 1954 1233 1958 1237
rect 484 1216 489 1219
rect 323 1193 328 1211
rect 341 1205 346 1211
rect 1872 1213 1877 1232
rect 406 1193 411 1211
rect 323 1188 411 1193
rect 424 1176 429 1211
rect 484 1202 489 1211
rect 1895 1213 1900 1232
rect 1953 1229 1958 1233
rect 2090 1233 2094 1237
rect 2236 1235 2240 1239
rect 1953 1219 1958 1224
rect 2008 1213 2013 1232
rect 2031 1213 2036 1232
rect 2089 1229 2094 1233
rect 2089 1219 2094 1224
rect 2154 1215 2159 1234
rect 2177 1215 2182 1234
rect 2235 1231 2240 1235
rect 2383 1235 2387 1239
rect 2513 1238 2518 1262
rect 2536 1238 2541 1262
rect 2594 1252 2599 1255
rect 2594 1238 2599 1247
rect 2649 1238 2654 1262
rect 2672 1238 2677 1262
rect 2730 1252 2735 1255
rect 2730 1238 2735 1247
rect 2795 1240 2800 1264
rect 2818 1240 2823 1264
rect 2876 1254 2881 1257
rect 2876 1240 2881 1249
rect 2942 1240 2947 1264
rect 2965 1240 2970 1264
rect 3023 1254 3028 1257
rect 3023 1240 3028 1249
rect 2235 1221 2240 1226
rect 2301 1215 2306 1234
rect 2324 1215 2329 1234
rect 2382 1231 2387 1235
rect 2595 1234 2599 1238
rect 2382 1221 2387 1226
rect 2513 1214 2518 1233
rect 2536 1214 2541 1233
rect 2594 1230 2599 1234
rect 2731 1234 2735 1238
rect 2877 1236 2881 1240
rect 2594 1220 2599 1225
rect 2649 1214 2654 1233
rect 2672 1214 2677 1233
rect 2730 1230 2735 1234
rect 2730 1220 2735 1225
rect 2795 1216 2800 1235
rect 2818 1216 2823 1235
rect 2876 1232 2881 1236
rect 3024 1236 3028 1240
rect 2876 1222 2881 1227
rect 2942 1216 2947 1235
rect 2965 1216 2970 1235
rect 3023 1232 3028 1236
rect 3023 1222 3028 1227
rect 485 1198 489 1202
rect 484 1194 489 1198
rect 484 1184 489 1189
rect 1872 1158 1877 1172
rect 1895 1158 1900 1172
rect 2016 1158 2021 1172
rect 2039 1158 2044 1172
rect 2165 1160 2170 1174
rect 2188 1160 2193 1174
rect 2310 1161 2315 1175
rect 2333 1161 2338 1175
rect 1872 1129 1877 1153
rect 1895 1129 1900 1153
rect 1953 1143 1958 1146
rect 1953 1129 1958 1138
rect 2016 1129 2021 1153
rect 2039 1129 2044 1153
rect 2097 1143 2102 1146
rect 2097 1129 2102 1138
rect 2165 1131 2170 1155
rect 2188 1131 2193 1155
rect 2246 1145 2251 1148
rect 2246 1131 2251 1140
rect 2310 1132 2315 1156
rect 2333 1132 2338 1156
rect 2391 1146 2396 1149
rect 2391 1132 2396 1141
rect 1954 1125 1958 1129
rect 1872 1105 1877 1124
rect 1565 1088 1570 1102
rect 1588 1088 1593 1102
rect 1895 1105 1900 1124
rect 1953 1121 1958 1125
rect 2098 1125 2102 1129
rect 2247 1127 2251 1131
rect 2392 1128 2396 1132
rect 1953 1111 1958 1116
rect 2016 1105 2021 1124
rect 2039 1105 2044 1124
rect 2097 1121 2102 1125
rect 2097 1111 2102 1116
rect 2165 1107 2170 1126
rect 2188 1107 2193 1126
rect 2246 1123 2251 1127
rect 2246 1113 2251 1118
rect 2310 1108 2315 1127
rect 2333 1108 2338 1127
rect 2391 1124 2396 1128
rect 2391 1114 2396 1119
rect 338 1054 376 1055
rect 381 1054 426 1055
rect 338 1050 426 1054
rect 209 1037 214 1040
rect 269 1037 274 1040
rect 320 1033 325 1037
rect 338 1033 343 1050
rect 403 1033 408 1037
rect 421 1033 426 1050
rect 751 1046 756 1060
rect 774 1046 779 1060
rect 898 1046 903 1060
rect 921 1046 926 1060
rect 1565 1059 1570 1083
rect 1588 1059 1593 1083
rect 1644 1074 1649 1077
rect 1644 1060 1649 1069
rect 1044 1044 1049 1058
rect 1067 1044 1072 1058
rect 1180 1044 1185 1058
rect 1203 1044 1208 1058
rect 1645 1056 1649 1060
rect 209 1023 214 1032
rect 210 1019 214 1023
rect 209 1015 214 1019
rect 269 1023 274 1032
rect 693 1031 698 1034
rect 269 1019 273 1023
rect 269 1015 274 1019
rect 320 1016 325 1028
rect 338 1024 343 1028
rect 403 1016 408 1028
rect 421 1024 426 1028
rect 693 1017 698 1026
rect 751 1017 756 1041
rect 774 1017 779 1041
rect 840 1031 845 1034
rect 840 1017 845 1026
rect 898 1017 903 1041
rect 921 1017 926 1041
rect 986 1029 991 1032
rect 321 1011 343 1016
rect 403 1011 426 1016
rect 209 1005 214 1010
rect 269 1005 274 1010
rect 301 999 325 1004
rect 301 991 306 999
rect 320 994 325 999
rect 338 994 343 1011
rect 403 994 408 998
rect 421 994 426 1011
rect 693 1013 697 1017
rect 693 1009 698 1013
rect 840 1013 844 1017
rect 693 999 698 1004
rect 481 994 486 997
rect 751 993 756 1012
rect 320 971 325 989
rect 338 983 343 989
rect 403 971 408 989
rect 320 966 408 971
rect 421 954 426 989
rect 481 980 486 989
rect 774 993 779 1012
rect 840 1009 845 1013
rect 986 1015 991 1024
rect 1044 1015 1049 1039
rect 1067 1015 1072 1039
rect 1122 1029 1127 1032
rect 1122 1015 1127 1024
rect 1180 1015 1185 1039
rect 1203 1015 1208 1039
rect 1565 1035 1570 1054
rect 1588 1035 1593 1054
rect 1644 1052 1649 1056
rect 1644 1043 1649 1047
rect 840 999 845 1004
rect 898 993 903 1012
rect 921 993 926 1012
rect 986 1011 990 1015
rect 986 1007 991 1011
rect 1122 1011 1126 1015
rect 986 997 991 1002
rect 1044 991 1049 1010
rect 1067 991 1072 1010
rect 1122 1007 1127 1011
rect 1122 997 1127 1002
rect 1180 991 1185 1010
rect 1203 991 1208 1010
rect 482 976 486 980
rect 481 972 486 976
rect 1564 970 1569 984
rect 1587 970 1592 984
rect 2273 978 2278 992
rect 2296 978 2301 992
rect 2409 978 2414 992
rect 2432 978 2437 992
rect 2555 980 2560 994
rect 2578 980 2583 994
rect 2702 980 2707 994
rect 2725 980 2730 994
rect 481 962 486 967
rect 742 939 747 953
rect 765 939 770 953
rect 887 938 892 952
rect 910 938 915 952
rect 684 924 689 927
rect 684 910 689 919
rect 742 910 747 934
rect 765 910 770 934
rect 1036 936 1041 950
rect 1059 936 1064 950
rect 1180 936 1185 950
rect 1203 936 1208 950
rect 1564 941 1569 965
rect 1587 941 1592 965
rect 1643 955 1648 958
rect 1643 941 1648 950
rect 2273 949 2278 973
rect 2296 949 2301 973
rect 2354 963 2359 966
rect 2354 949 2359 958
rect 2409 949 2414 973
rect 2432 949 2437 973
rect 2490 963 2495 966
rect 2490 949 2495 958
rect 2555 951 2560 975
rect 2578 951 2583 975
rect 2636 965 2641 968
rect 2636 951 2641 960
rect 2702 951 2707 975
rect 2725 951 2730 975
rect 2783 965 2788 968
rect 2783 951 2788 960
rect 2355 945 2359 949
rect 829 923 834 926
rect 684 906 688 910
rect 684 902 689 906
rect 829 909 834 918
rect 887 909 892 933
rect 910 909 915 933
rect 1416 935 1421 938
rect 1454 935 1459 938
rect 1644 937 1648 941
rect 978 921 983 924
rect 829 905 833 909
rect 684 892 689 897
rect 742 886 747 905
rect 765 886 770 905
rect 829 901 834 905
rect 978 907 983 916
rect 1036 907 1041 931
rect 1059 907 1064 931
rect 1122 921 1127 924
rect 1122 907 1127 916
rect 1180 907 1185 931
rect 1203 907 1208 931
rect 1416 921 1421 930
rect 1454 921 1459 930
rect 1417 917 1421 921
rect 1455 917 1459 921
rect 1416 913 1421 917
rect 1454 913 1459 917
rect 1564 917 1569 936
rect 1587 917 1592 936
rect 1643 933 1648 937
rect 1643 923 1648 928
rect 829 891 834 896
rect 887 885 892 904
rect 910 885 915 904
rect 978 903 982 907
rect 978 899 983 903
rect 1122 903 1126 907
rect 978 889 983 894
rect 1036 883 1041 902
rect 18 864 23 867
rect 77 860 82 879
rect 93 860 98 879
rect 1059 883 1064 902
rect 1122 899 1127 903
rect 1416 903 1421 908
rect 1454 903 1459 908
rect 1122 889 1127 894
rect 1180 883 1185 902
rect 1203 883 1208 902
rect 2012 900 2017 908
rect 2036 900 2041 934
rect 2273 925 2278 944
rect 2296 925 2301 944
rect 2354 941 2359 945
rect 2491 945 2495 949
rect 2637 947 2641 951
rect 2354 931 2359 936
rect 2409 925 2414 944
rect 2432 925 2437 944
rect 2490 941 2495 945
rect 2490 931 2495 936
rect 2555 927 2560 946
rect 2578 927 2583 946
rect 2636 943 2641 947
rect 2784 947 2788 951
rect 2636 933 2641 938
rect 2702 927 2707 946
rect 2725 927 2730 946
rect 2783 943 2788 947
rect 2783 933 2788 938
rect 2081 902 2086 905
rect 2012 885 2017 895
rect 2013 880 2017 885
rect 341 869 379 870
rect 384 869 429 870
rect 341 865 429 869
rect 1563 866 1568 880
rect 1586 866 1591 880
rect 109 860 114 864
rect 125 860 130 864
rect 18 850 23 859
rect 18 846 22 850
rect 18 842 23 846
rect 18 832 23 837
rect 77 826 82 855
rect 93 826 98 855
rect 109 826 114 855
rect 125 826 130 855
rect 212 852 217 855
rect 272 852 277 855
rect 323 848 328 852
rect 341 848 346 865
rect 406 848 411 852
rect 424 848 429 865
rect 2012 863 2017 880
rect 2036 863 2041 895
rect 2081 888 2086 897
rect 2082 884 2086 888
rect 2081 880 2086 884
rect 2081 870 2086 875
rect 2273 870 2278 884
rect 2296 870 2301 884
rect 2417 870 2422 884
rect 2440 870 2445 884
rect 2566 872 2571 886
rect 2589 872 2594 886
rect 2711 873 2716 887
rect 2734 873 2739 887
rect 212 838 217 847
rect 213 834 217 838
rect 212 830 217 834
rect 272 838 277 847
rect 272 834 276 838
rect 272 830 277 834
rect 323 831 328 843
rect 341 839 346 843
rect 406 831 411 843
rect 424 839 429 843
rect 1563 837 1568 861
rect 1586 837 1591 861
rect 2012 854 2017 858
rect 2036 854 2041 858
rect 1644 851 1649 854
rect 1644 837 1649 846
rect 2273 841 2278 865
rect 2296 841 2301 865
rect 2354 855 2359 858
rect 2354 841 2359 850
rect 2417 841 2422 865
rect 2440 841 2445 865
rect 2498 855 2503 858
rect 2498 841 2503 850
rect 2566 843 2571 867
rect 2589 843 2594 867
rect 2647 857 2652 860
rect 2647 843 2652 852
rect 2711 844 2716 868
rect 2734 844 2739 868
rect 2792 858 2797 861
rect 2792 844 2797 853
rect 1645 833 1649 837
rect 2355 837 2359 841
rect 324 826 346 831
rect 406 826 429 831
rect 77 814 82 821
rect 93 814 98 821
rect 109 804 114 821
rect 125 804 130 821
rect 212 820 217 825
rect 272 820 277 825
rect 304 814 328 819
rect 304 806 309 814
rect 323 809 328 814
rect 341 809 346 826
rect 406 809 411 813
rect 424 809 429 826
rect 1563 813 1568 832
rect 484 809 489 812
rect 323 786 328 804
rect 341 798 346 804
rect 1586 813 1591 832
rect 1644 829 1649 833
rect 1644 819 1649 824
rect 2273 817 2278 836
rect 2296 817 2301 836
rect 2354 833 2359 837
rect 2499 837 2503 841
rect 2648 839 2652 843
rect 2793 840 2797 844
rect 2354 823 2359 828
rect 2417 817 2422 836
rect 2440 817 2445 836
rect 2498 833 2503 837
rect 2498 823 2503 828
rect 2566 819 2571 838
rect 2589 819 2594 838
rect 2647 835 2652 839
rect 2647 825 2652 830
rect 2711 820 2716 839
rect 2734 820 2739 839
rect 2792 836 2797 840
rect 2792 826 2797 831
rect 406 786 411 804
rect 323 781 411 786
rect 424 769 429 804
rect 484 795 489 804
rect 485 791 489 795
rect 484 787 489 791
rect 484 777 489 782
rect 1563 770 1568 784
rect 1586 770 1591 784
rect 1563 741 1568 765
rect 1586 741 1591 765
rect 1643 755 1648 758
rect 1643 741 1648 750
rect 1644 737 1648 741
rect 1563 717 1568 736
rect 1586 717 1591 736
rect 1643 733 1648 737
rect 1643 723 1648 728
rect 341 694 379 695
rect 384 694 429 695
rect 341 690 429 694
rect 212 677 217 680
rect 272 677 277 680
rect 323 673 328 677
rect 341 673 346 690
rect 406 673 411 677
rect 424 673 429 690
rect 212 663 217 672
rect 213 659 217 663
rect 212 655 217 659
rect 272 663 277 672
rect 272 659 276 663
rect 272 655 277 659
rect 323 656 328 668
rect 341 664 346 668
rect 406 656 411 668
rect 424 664 429 668
rect 2097 664 2135 665
rect 2140 664 2185 665
rect 2097 660 2185 664
rect 324 651 346 656
rect 406 651 429 656
rect 212 645 217 650
rect 272 645 277 650
rect 304 639 328 644
rect 304 631 309 639
rect 323 634 328 639
rect 341 634 346 651
rect 406 634 411 638
rect 424 634 429 651
rect 2024 647 2029 650
rect 2079 643 2084 647
rect 2097 643 2102 660
rect 2162 643 2167 647
rect 2180 643 2185 660
rect 484 634 489 637
rect 2024 633 2029 642
rect 2024 629 2028 633
rect 323 611 328 629
rect 341 623 346 629
rect 406 611 411 629
rect 323 606 411 611
rect 424 594 429 629
rect 484 620 489 629
rect 2024 625 2029 629
rect 2079 626 2084 638
rect 2097 634 2102 638
rect 2162 626 2167 638
rect 2180 634 2185 638
rect 2080 621 2102 626
rect 2162 621 2185 626
rect 485 616 489 620
rect 484 612 489 616
rect 2024 615 2029 620
rect 2060 609 2084 614
rect 484 602 489 607
rect 2060 601 2065 609
rect 2079 604 2084 609
rect 2097 604 2102 621
rect 2162 604 2167 608
rect 2180 604 2185 621
rect 2240 604 2245 607
rect 2079 581 2084 599
rect 2097 593 2102 599
rect 2162 581 2167 599
rect 2079 576 2167 581
rect 2180 564 2185 599
rect 2240 590 2245 599
rect 2241 586 2245 590
rect 2240 582 2245 586
rect 2240 572 2245 577
rect 1476 541 1481 544
rect 1539 537 1544 540
rect 1555 537 1560 540
rect 1571 537 1576 540
rect 1476 527 1481 536
rect 1476 523 1480 527
rect 1476 519 1481 523
rect 1476 509 1481 514
rect 1539 501 1544 532
rect 1555 501 1560 532
rect 1571 501 1576 532
rect 1539 485 1544 496
rect 1555 485 1560 496
rect 1571 485 1576 496
rect 2091 481 2129 482
rect 2134 481 2179 482
rect 2091 477 2179 481
rect 2018 464 2023 467
rect 2073 460 2078 464
rect 2091 460 2096 477
rect 2156 460 2161 464
rect 2174 460 2179 477
rect 2018 450 2023 459
rect 2018 446 2022 450
rect 2018 442 2023 446
rect 2073 443 2078 455
rect 2091 451 2096 455
rect 2156 443 2161 455
rect 2174 451 2179 455
rect 2074 438 2096 443
rect 2156 438 2179 443
rect 1360 423 1365 437
rect 1383 423 1388 437
rect 1506 421 1511 435
rect 1529 421 1534 435
rect 1642 421 1647 435
rect 1665 421 1670 435
rect 2018 432 2023 437
rect 2054 426 2078 431
rect 1302 408 1307 411
rect 1302 394 1307 403
rect 1360 394 1365 418
rect 1383 394 1388 418
rect 2054 418 2059 426
rect 2073 421 2078 426
rect 2091 421 2096 438
rect 2156 421 2161 425
rect 2174 421 2179 438
rect 2234 421 2239 424
rect 1448 406 1453 409
rect 1302 390 1306 394
rect 1302 386 1307 390
rect 1448 392 1453 401
rect 1506 392 1511 416
rect 1529 392 1534 416
rect 1584 406 1589 409
rect 1584 392 1589 401
rect 1642 392 1647 416
rect 1665 392 1670 416
rect 2073 398 2078 416
rect 2091 410 2096 416
rect 2156 398 2161 416
rect 2073 393 2161 398
rect 1302 376 1307 381
rect 1360 370 1365 389
rect 1383 370 1388 389
rect 1448 388 1452 392
rect 1448 384 1453 388
rect 1584 388 1588 392
rect 1448 374 1453 379
rect 1506 368 1511 387
rect 1529 368 1534 387
rect 1584 384 1589 388
rect 1584 374 1589 379
rect 1642 368 1647 387
rect 1665 368 1670 387
rect 2174 381 2179 416
rect 2234 407 2239 416
rect 2235 403 2239 407
rect 2234 399 2239 403
rect 2234 389 2239 394
rect 2079 309 2117 310
rect 2122 309 2167 310
rect 2079 305 2167 309
rect 1310 292 1355 293
rect 1360 292 1398 293
rect 1310 288 1398 292
rect 1310 271 1315 288
rect 1328 271 1333 275
rect 1393 271 1398 288
rect 1648 292 1693 293
rect 1698 292 1736 293
rect 2006 292 2011 295
rect 1648 288 1736 292
rect 1474 275 1479 278
rect 1411 271 1416 275
rect 1648 271 1653 288
rect 1666 271 1671 275
rect 1731 271 1736 288
rect 2061 288 2066 292
rect 2079 288 2084 305
rect 2144 288 2149 292
rect 2162 288 2167 305
rect 2006 278 2011 287
rect 1806 275 1811 278
rect 1749 271 1754 275
rect 1310 262 1315 266
rect 1328 254 1333 266
rect 1393 262 1398 266
rect 1411 254 1416 266
rect 1474 261 1479 270
rect 2006 274 2010 278
rect 2006 270 2011 274
rect 2061 271 2066 283
rect 2079 279 2084 283
rect 2144 271 2149 283
rect 2162 279 2167 283
rect 1648 262 1653 266
rect 1475 257 1479 261
rect 1310 249 1333 254
rect 1393 249 1415 254
rect 1474 253 1479 257
rect 1666 254 1671 266
rect 1731 262 1736 266
rect 1749 254 1754 266
rect 1806 261 1811 270
rect 2062 266 2084 271
rect 2144 266 2167 271
rect 1807 257 1811 261
rect 2006 260 2011 265
rect 1250 232 1255 235
rect 1310 232 1315 249
rect 1328 232 1333 236
rect 1393 232 1398 249
rect 1648 249 1671 254
rect 1731 249 1753 254
rect 1806 253 1811 257
rect 2042 254 2066 259
rect 1474 243 1479 248
rect 1411 237 1435 242
rect 1411 232 1416 237
rect 1430 229 1435 237
rect 1588 232 1593 235
rect 1648 232 1653 249
rect 1666 232 1671 236
rect 1731 232 1736 249
rect 1806 243 1811 248
rect 2042 246 2047 254
rect 2061 249 2066 254
rect 2079 249 2084 266
rect 2144 249 2149 253
rect 2162 249 2167 266
rect 2222 249 2227 252
rect 1749 237 1773 242
rect 1749 232 1754 237
rect 1250 218 1255 227
rect 1250 214 1254 218
rect 1250 210 1255 214
rect 1250 200 1255 205
rect 1310 192 1315 227
rect 1328 209 1333 227
rect 1393 221 1398 227
rect 1411 209 1416 227
rect 1588 218 1593 227
rect 1588 214 1592 218
rect 1588 210 1593 214
rect 1328 204 1416 209
rect 1588 200 1593 205
rect 1648 192 1653 227
rect 1666 209 1671 227
rect 1768 229 1773 237
rect 1731 221 1736 227
rect 1749 209 1754 227
rect 2061 226 2066 244
rect 2079 238 2084 244
rect 2144 226 2149 244
rect 2061 221 2149 226
rect 1666 204 1754 209
rect 2162 209 2167 244
rect 2222 235 2227 244
rect 2223 231 2227 235
rect 2222 227 2227 231
rect 2222 217 2227 222
rect 2070 125 2108 126
rect 2113 125 2158 126
rect 2070 121 2158 125
rect 1997 108 2002 111
rect 2052 104 2057 108
rect 2070 104 2075 121
rect 2135 104 2140 108
rect 2153 104 2158 121
rect 1997 94 2002 103
rect 1997 90 2001 94
rect 1997 86 2002 90
rect 2052 87 2057 99
rect 2070 95 2075 99
rect 2135 87 2140 99
rect 2153 95 2158 99
rect 2053 82 2075 87
rect 2135 82 2158 87
rect 1997 76 2002 81
rect 2033 70 2057 75
rect 2033 62 2038 70
rect 2052 65 2057 70
rect 2070 65 2075 82
rect 2135 65 2140 69
rect 2153 65 2158 82
rect 2213 65 2218 68
rect 2052 42 2057 60
rect 2070 54 2075 60
rect 2135 42 2140 60
rect 2052 37 2140 42
rect 2153 25 2158 60
rect 2213 51 2218 60
rect 2214 47 2218 51
rect 2213 43 2218 47
rect 2213 33 2218 38
rect 1444 20 1449 23
rect 1507 16 1512 19
rect 1523 16 1528 19
rect 1539 16 1544 19
rect 1444 6 1449 15
rect 1444 2 1448 6
rect 1444 -2 1449 2
rect 1444 -12 1449 -7
rect 1507 -20 1512 11
rect 1523 -20 1528 11
rect 1539 -20 1544 11
rect 1507 -36 1512 -25
rect 1523 -36 1528 -25
rect 1539 -36 1544 -25
rect 1328 -98 1333 -84
rect 1351 -98 1356 -84
rect 1474 -100 1479 -86
rect 1497 -100 1502 -86
rect 1610 -100 1615 -86
rect 1633 -100 1638 -86
rect 1270 -113 1275 -110
rect 1270 -127 1275 -118
rect 1328 -127 1333 -103
rect 1351 -127 1356 -103
rect 1416 -115 1421 -112
rect 1270 -131 1274 -127
rect 1270 -135 1275 -131
rect 1416 -129 1421 -120
rect 1474 -129 1479 -105
rect 1497 -129 1502 -105
rect 1552 -115 1557 -112
rect 1552 -129 1557 -120
rect 1610 -129 1615 -105
rect 1633 -129 1638 -105
rect 1270 -145 1275 -140
rect 1328 -151 1333 -132
rect 1351 -151 1356 -132
rect 1416 -133 1420 -129
rect 1416 -137 1421 -133
rect 1552 -133 1556 -129
rect 1416 -147 1421 -142
rect 1474 -153 1479 -134
rect 1497 -153 1502 -134
rect 1552 -137 1557 -133
rect 1552 -147 1557 -142
rect 1610 -153 1615 -134
rect 1633 -153 1638 -134
rect 1278 -229 1323 -228
rect 1328 -229 1366 -228
rect 1278 -233 1366 -229
rect 1278 -250 1283 -233
rect 1296 -250 1301 -246
rect 1361 -250 1366 -233
rect 1616 -229 1661 -228
rect 1666 -229 1704 -228
rect 1616 -233 1704 -229
rect 1442 -246 1447 -243
rect 1379 -250 1384 -246
rect 1616 -250 1621 -233
rect 1634 -250 1639 -246
rect 1699 -250 1704 -233
rect 1774 -246 1779 -243
rect 1717 -250 1722 -246
rect 1278 -259 1283 -255
rect 1296 -267 1301 -255
rect 1361 -259 1366 -255
rect 1379 -267 1384 -255
rect 1442 -260 1447 -251
rect 1616 -259 1621 -255
rect 1443 -264 1447 -260
rect 1278 -272 1301 -267
rect 1361 -272 1383 -267
rect 1442 -268 1447 -264
rect 1634 -267 1639 -255
rect 1699 -259 1704 -255
rect 1717 -267 1722 -255
rect 1774 -260 1779 -251
rect 1775 -264 1779 -260
rect 1218 -289 1223 -286
rect 1278 -289 1283 -272
rect 1296 -289 1301 -285
rect 1361 -289 1366 -272
rect 1616 -272 1639 -267
rect 1699 -272 1721 -267
rect 1774 -268 1779 -264
rect 1442 -278 1447 -273
rect 1379 -284 1403 -279
rect 1379 -289 1384 -284
rect 1218 -303 1223 -294
rect 1218 -307 1222 -303
rect 1218 -311 1223 -307
rect 1218 -321 1223 -316
rect 1278 -329 1283 -294
rect 1296 -312 1301 -294
rect 1398 -292 1403 -284
rect 1556 -289 1561 -286
rect 1616 -289 1621 -272
rect 1634 -289 1639 -285
rect 1699 -289 1704 -272
rect 1774 -278 1779 -273
rect 1717 -284 1741 -279
rect 1717 -289 1722 -284
rect 1361 -300 1366 -294
rect 1379 -312 1384 -294
rect 1556 -303 1561 -294
rect 1556 -307 1560 -303
rect 1556 -311 1561 -307
rect 1296 -317 1384 -312
rect 1556 -321 1561 -316
rect 1616 -329 1621 -294
rect 1634 -312 1639 -294
rect 1736 -292 1741 -284
rect 1699 -300 1704 -294
rect 1717 -312 1722 -294
rect 1634 -317 1722 -312
rect 1444 -431 1449 -428
rect 1507 -435 1512 -432
rect 1523 -435 1528 -432
rect 1539 -435 1544 -432
rect 1444 -445 1449 -436
rect 1444 -449 1448 -445
rect 1444 -453 1449 -449
rect 1444 -463 1449 -458
rect 1507 -471 1512 -440
rect 1523 -471 1528 -440
rect 1539 -471 1544 -440
rect 1507 -487 1512 -476
rect 1523 -487 1528 -476
rect 1539 -487 1544 -476
rect 1328 -549 1333 -535
rect 1351 -549 1356 -535
rect 1474 -551 1479 -537
rect 1497 -551 1502 -537
rect 1610 -551 1615 -537
rect 1633 -551 1638 -537
rect 1270 -564 1275 -561
rect 1270 -578 1275 -569
rect 1328 -578 1333 -554
rect 1351 -578 1356 -554
rect 1416 -566 1421 -563
rect 1270 -582 1274 -578
rect 1270 -586 1275 -582
rect 1416 -580 1421 -571
rect 1474 -580 1479 -556
rect 1497 -580 1502 -556
rect 1552 -566 1557 -563
rect 1552 -580 1557 -571
rect 1610 -580 1615 -556
rect 1633 -580 1638 -556
rect 1270 -596 1275 -591
rect 1328 -602 1333 -583
rect 1351 -602 1356 -583
rect 1416 -584 1420 -580
rect 1416 -588 1421 -584
rect 1552 -584 1556 -580
rect 1416 -598 1421 -593
rect 1474 -604 1479 -585
rect 1497 -604 1502 -585
rect 1552 -588 1557 -584
rect 1552 -598 1557 -593
rect 1610 -604 1615 -585
rect 1633 -604 1638 -585
rect 1278 -680 1323 -679
rect 1328 -680 1366 -679
rect 1278 -684 1366 -680
rect 1278 -701 1283 -684
rect 1296 -701 1301 -697
rect 1361 -701 1366 -684
rect 1616 -680 1661 -679
rect 1666 -680 1704 -679
rect 1616 -684 1704 -680
rect 1442 -697 1447 -694
rect 1379 -701 1384 -697
rect 1616 -701 1621 -684
rect 1634 -701 1639 -697
rect 1699 -701 1704 -684
rect 1774 -697 1779 -694
rect 1717 -701 1722 -697
rect 1278 -710 1283 -706
rect 1296 -718 1301 -706
rect 1361 -710 1366 -706
rect 1379 -718 1384 -706
rect 1442 -711 1447 -702
rect 1616 -710 1621 -706
rect 1443 -715 1447 -711
rect 1278 -723 1301 -718
rect 1361 -723 1383 -718
rect 1442 -719 1447 -715
rect 1634 -718 1639 -706
rect 1699 -710 1704 -706
rect 1717 -718 1722 -706
rect 1774 -711 1779 -702
rect 1775 -715 1779 -711
rect 1218 -740 1223 -737
rect 1278 -740 1283 -723
rect 1296 -740 1301 -736
rect 1361 -740 1366 -723
rect 1616 -723 1639 -718
rect 1699 -723 1721 -718
rect 1774 -719 1779 -715
rect 1442 -729 1447 -724
rect 1379 -735 1403 -730
rect 1379 -740 1384 -735
rect 1218 -754 1223 -745
rect 1218 -758 1222 -754
rect 1218 -762 1223 -758
rect 1218 -772 1223 -767
rect 1278 -780 1283 -745
rect 1296 -763 1301 -745
rect 1398 -743 1403 -735
rect 1556 -740 1561 -737
rect 1616 -740 1621 -723
rect 1634 -740 1639 -736
rect 1361 -751 1366 -745
rect 1379 -763 1384 -745
rect 1699 -740 1704 -723
rect 1774 -729 1779 -724
rect 1717 -735 1741 -730
rect 1717 -740 1722 -735
rect 1736 -743 1741 -735
rect 1556 -754 1561 -745
rect 1556 -758 1560 -754
rect 1556 -762 1561 -758
rect 1296 -768 1384 -763
rect 1556 -772 1561 -767
rect 1616 -780 1621 -745
rect 1634 -763 1639 -745
rect 1699 -751 1704 -745
rect 1717 -763 1722 -745
rect 1634 -768 1722 -763
rect 1435 -881 1440 -878
rect 1498 -885 1503 -882
rect 1514 -885 1519 -882
rect 1530 -885 1535 -882
rect 1435 -895 1440 -886
rect 1435 -899 1439 -895
rect 1435 -903 1440 -899
rect 1435 -913 1440 -908
rect 1498 -921 1503 -890
rect 1514 -921 1519 -890
rect 1530 -921 1535 -890
rect 1498 -937 1503 -926
rect 1514 -937 1519 -926
rect 1530 -937 1535 -926
rect 1319 -999 1324 -985
rect 1342 -999 1347 -985
rect 1465 -1001 1470 -987
rect 1488 -1001 1493 -987
rect 1601 -1001 1606 -987
rect 1624 -1001 1629 -987
rect 1261 -1014 1266 -1011
rect 1261 -1028 1266 -1019
rect 1319 -1028 1324 -1004
rect 1342 -1028 1347 -1004
rect 1407 -1016 1412 -1013
rect 1261 -1032 1265 -1028
rect 1261 -1036 1266 -1032
rect 1407 -1030 1412 -1021
rect 1465 -1030 1470 -1006
rect 1488 -1030 1493 -1006
rect 1543 -1016 1548 -1013
rect 1543 -1030 1548 -1021
rect 1601 -1030 1606 -1006
rect 1624 -1030 1629 -1006
rect 1261 -1046 1266 -1041
rect 1319 -1052 1324 -1033
rect 1342 -1052 1347 -1033
rect 1407 -1034 1411 -1030
rect 1407 -1038 1412 -1034
rect 1543 -1034 1547 -1030
rect 1407 -1048 1412 -1043
rect 1465 -1054 1470 -1035
rect 1488 -1054 1493 -1035
rect 1543 -1038 1548 -1034
rect 1543 -1048 1548 -1043
rect 1601 -1054 1606 -1035
rect 1624 -1054 1629 -1035
rect 1269 -1130 1314 -1129
rect 1319 -1130 1357 -1129
rect 1269 -1134 1357 -1130
rect 1269 -1151 1274 -1134
rect 1287 -1151 1292 -1147
rect 1352 -1151 1357 -1134
rect 1607 -1130 1652 -1129
rect 1657 -1130 1695 -1129
rect 1607 -1134 1695 -1130
rect 1433 -1147 1438 -1144
rect 1370 -1151 1375 -1147
rect 1607 -1151 1612 -1134
rect 1625 -1151 1630 -1147
rect 1690 -1151 1695 -1134
rect 1765 -1147 1770 -1144
rect 1708 -1151 1713 -1147
rect 1269 -1160 1274 -1156
rect 1287 -1168 1292 -1156
rect 1352 -1160 1357 -1156
rect 1370 -1168 1375 -1156
rect 1433 -1161 1438 -1152
rect 1607 -1160 1612 -1156
rect 1434 -1165 1438 -1161
rect 1269 -1173 1292 -1168
rect 1352 -1173 1374 -1168
rect 1433 -1169 1438 -1165
rect 1625 -1168 1630 -1156
rect 1690 -1160 1695 -1156
rect 1708 -1168 1713 -1156
rect 1765 -1161 1770 -1152
rect 1766 -1165 1770 -1161
rect 1209 -1190 1214 -1187
rect 1269 -1190 1274 -1173
rect 1287 -1190 1292 -1186
rect 1352 -1190 1357 -1173
rect 1607 -1173 1630 -1168
rect 1690 -1173 1712 -1168
rect 1765 -1169 1770 -1165
rect 1433 -1179 1438 -1174
rect 1370 -1185 1394 -1180
rect 1370 -1190 1375 -1185
rect 1389 -1193 1394 -1185
rect 1547 -1190 1552 -1187
rect 1607 -1190 1612 -1173
rect 1625 -1190 1630 -1186
rect 1690 -1190 1695 -1173
rect 1765 -1179 1770 -1174
rect 1708 -1185 1732 -1180
rect 1708 -1190 1713 -1185
rect 1209 -1204 1214 -1195
rect 1209 -1208 1213 -1204
rect 1209 -1212 1214 -1208
rect 1209 -1222 1214 -1217
rect 1269 -1230 1274 -1195
rect 1287 -1213 1292 -1195
rect 1352 -1201 1357 -1195
rect 1370 -1213 1375 -1195
rect 1547 -1204 1552 -1195
rect 1547 -1208 1551 -1204
rect 1547 -1212 1552 -1208
rect 1287 -1218 1375 -1213
rect 1547 -1222 1552 -1217
rect 1607 -1230 1612 -1195
rect 1625 -1213 1630 -1195
rect 1727 -1193 1732 -1185
rect 1690 -1201 1695 -1195
rect 1708 -1213 1713 -1195
rect 1625 -1218 1713 -1213
<< polycontact >>
rect 882 1562 887 1566
rect 936 1536 941 1542
rect 959 1536 964 1542
rect 774 1480 779 1484
rect 831 1481 836 1485
rect 669 1435 674 1442
rect 685 1435 690 1442
rect 701 1435 706 1442
rect 717 1436 722 1443
rect 722 1310 727 1315
rect 738 1310 744 1316
rect 883 1310 889 1317
rect 899 1310 905 1317
rect 931 1310 937 1316
rect 1060 1312 1067 1318
rect 379 1276 384 1281
rect 639 1277 644 1281
rect 1075 1310 1085 1318
rect 828 1277 833 1281
rect 986 1277 991 1281
rect 208 1241 213 1245
rect 1144 1259 1149 1263
rect 276 1241 281 1245
rect 319 1233 324 1238
rect 915 1229 922 1235
rect 1043 1229 1051 1236
rect 1198 1233 1203 1239
rect 1221 1233 1226 1239
rect 1949 1233 1954 1237
rect 304 1208 309 1213
rect 1872 1207 1877 1213
rect 2085 1233 2090 1237
rect 2231 1235 2236 1239
rect 1895 1207 1900 1213
rect 2008 1207 2013 1213
rect 2031 1207 2036 1213
rect 2154 1209 2159 1215
rect 2378 1235 2383 1239
rect 2177 1209 2182 1215
rect 2301 1209 2306 1215
rect 2590 1234 2595 1238
rect 2324 1209 2329 1215
rect 2513 1208 2518 1214
rect 2726 1234 2731 1238
rect 2872 1236 2877 1240
rect 2536 1208 2541 1214
rect 2649 1208 2654 1214
rect 2672 1208 2677 1214
rect 2795 1210 2800 1216
rect 3019 1236 3024 1240
rect 2818 1210 2823 1216
rect 2942 1210 2947 1216
rect 2965 1210 2970 1216
rect 480 1198 485 1202
rect 424 1171 429 1176
rect 1949 1125 1954 1129
rect 1872 1099 1877 1105
rect 2093 1125 2098 1129
rect 2242 1127 2247 1131
rect 2387 1128 2392 1132
rect 1895 1099 1900 1105
rect 2016 1099 2021 1105
rect 2039 1099 2044 1105
rect 2165 1101 2170 1107
rect 2188 1101 2193 1107
rect 2310 1102 2315 1108
rect 2333 1102 2338 1108
rect 376 1054 381 1059
rect 1640 1056 1645 1060
rect 205 1019 210 1023
rect 273 1019 278 1023
rect 316 1011 321 1016
rect 301 986 306 991
rect 697 1013 702 1017
rect 844 1013 849 1017
rect 751 987 756 993
rect 1565 1029 1570 1035
rect 1588 1029 1593 1035
rect 774 987 779 993
rect 898 987 903 993
rect 990 1011 995 1015
rect 1126 1011 1131 1015
rect 921 987 926 993
rect 1044 985 1049 991
rect 1067 985 1072 991
rect 1180 985 1185 991
rect 1203 985 1208 991
rect 477 976 482 980
rect 421 949 426 954
rect 2350 945 2355 949
rect 688 906 693 910
rect 1639 937 1644 941
rect 833 905 838 909
rect 77 879 83 886
rect 93 879 99 886
rect 742 880 747 886
rect 1412 917 1417 921
rect 1450 917 1455 921
rect 1564 911 1569 917
rect 2036 934 2042 940
rect 1587 911 1592 917
rect 765 880 770 886
rect 887 879 892 885
rect 982 903 987 907
rect 1126 903 1131 907
rect 910 879 915 885
rect 1036 877 1041 883
rect 1059 877 1064 883
rect 1180 877 1185 883
rect 2273 919 2278 925
rect 2486 945 2491 949
rect 2632 947 2637 951
rect 2296 919 2301 925
rect 2409 919 2414 925
rect 2432 919 2437 925
rect 2555 921 2560 927
rect 2779 947 2784 951
rect 2578 921 2583 927
rect 2702 921 2707 927
rect 2725 921 2730 927
rect 1203 877 1208 883
rect 2008 880 2013 885
rect 379 869 384 874
rect 22 846 27 850
rect 2077 884 2082 888
rect 208 834 213 838
rect 276 834 281 838
rect 1640 833 1645 837
rect 2350 837 2355 841
rect 319 826 324 831
rect 109 798 116 804
rect 125 798 132 804
rect 304 801 309 806
rect 1563 807 1568 813
rect 1586 807 1591 813
rect 2273 811 2278 817
rect 2494 837 2499 841
rect 2643 839 2648 843
rect 2788 840 2793 844
rect 2296 811 2301 817
rect 2417 811 2422 817
rect 2440 811 2445 817
rect 2566 813 2571 819
rect 2589 813 2594 819
rect 2711 814 2716 820
rect 2734 814 2739 820
rect 480 791 485 795
rect 424 764 429 769
rect 1639 737 1644 741
rect 1563 711 1568 717
rect 1586 711 1591 717
rect 379 694 384 699
rect 208 659 213 663
rect 276 659 281 663
rect 2135 664 2140 669
rect 319 651 324 656
rect 304 626 309 631
rect 2028 629 2033 633
rect 2075 621 2080 626
rect 480 616 485 620
rect 2060 596 2065 601
rect 424 589 429 594
rect 2236 586 2241 590
rect 2180 559 2185 564
rect 1480 523 1485 527
rect 1539 478 1544 485
rect 1555 478 1560 485
rect 1571 478 1576 485
rect 2129 481 2134 486
rect 2022 446 2027 450
rect 2069 438 2074 443
rect 1306 390 1311 394
rect 2054 413 2059 418
rect 1360 364 1365 370
rect 1452 388 1457 392
rect 1588 388 1593 392
rect 1383 364 1388 370
rect 1506 362 1511 368
rect 1529 362 1534 368
rect 1642 362 1647 368
rect 2230 403 2235 407
rect 2174 376 2179 381
rect 1665 362 1670 368
rect 2117 309 2122 314
rect 1355 292 1360 297
rect 1693 292 1698 297
rect 2010 274 2015 278
rect 1470 257 1475 261
rect 1415 249 1420 254
rect 2057 266 2062 271
rect 1802 257 1807 261
rect 1753 249 1758 254
rect 2042 241 2047 246
rect 1254 214 1259 218
rect 1430 224 1435 229
rect 1592 214 1597 218
rect 1310 187 1315 192
rect 1768 224 1773 229
rect 2218 231 2223 235
rect 2162 204 2167 209
rect 1648 187 1653 192
rect 2108 125 2113 130
rect 2001 90 2006 94
rect 2048 82 2053 87
rect 2033 57 2038 62
rect 2209 47 2214 51
rect 2153 20 2158 25
rect 1448 2 1453 6
rect 1507 -43 1512 -36
rect 1523 -43 1528 -36
rect 1539 -43 1544 -36
rect 1274 -131 1279 -127
rect 1328 -157 1333 -151
rect 1420 -133 1425 -129
rect 1556 -133 1561 -129
rect 1351 -157 1356 -151
rect 1474 -159 1479 -153
rect 1497 -159 1502 -153
rect 1610 -159 1615 -153
rect 1633 -159 1638 -153
rect 1323 -229 1328 -224
rect 1661 -229 1666 -224
rect 1438 -264 1443 -260
rect 1383 -272 1388 -267
rect 1770 -264 1775 -260
rect 1721 -272 1726 -267
rect 1222 -307 1227 -303
rect 1398 -297 1403 -292
rect 1560 -307 1565 -303
rect 1278 -334 1283 -329
rect 1736 -297 1741 -292
rect 1616 -334 1621 -329
rect 1448 -449 1453 -445
rect 1507 -494 1512 -487
rect 1523 -494 1528 -487
rect 1539 -494 1544 -487
rect 1274 -582 1279 -578
rect 1328 -608 1333 -602
rect 1420 -584 1425 -580
rect 1556 -584 1561 -580
rect 1351 -608 1356 -602
rect 1474 -610 1479 -604
rect 1497 -610 1502 -604
rect 1610 -610 1615 -604
rect 1633 -610 1638 -604
rect 1323 -680 1328 -675
rect 1661 -680 1666 -675
rect 1438 -715 1443 -711
rect 1383 -723 1388 -718
rect 1770 -715 1775 -711
rect 1721 -723 1726 -718
rect 1222 -758 1227 -754
rect 1398 -748 1403 -743
rect 1560 -758 1565 -754
rect 1278 -785 1283 -780
rect 1736 -748 1741 -743
rect 1616 -785 1621 -780
rect 1439 -899 1444 -895
rect 1498 -944 1503 -937
rect 1514 -944 1519 -937
rect 1530 -944 1535 -937
rect 1265 -1032 1270 -1028
rect 1319 -1058 1324 -1052
rect 1411 -1034 1416 -1030
rect 1547 -1034 1552 -1030
rect 1342 -1058 1347 -1052
rect 1465 -1060 1470 -1054
rect 1488 -1060 1493 -1054
rect 1601 -1060 1606 -1054
rect 1624 -1060 1629 -1054
rect 1314 -1130 1319 -1125
rect 1652 -1130 1657 -1125
rect 1429 -1165 1434 -1161
rect 1374 -1173 1379 -1168
rect 1761 -1165 1766 -1161
rect 1712 -1173 1717 -1168
rect 1213 -1208 1218 -1204
rect 1389 -1198 1394 -1193
rect 1551 -1208 1556 -1204
rect 1269 -1235 1274 -1230
rect 1727 -1198 1732 -1193
rect 1607 -1235 1612 -1230
<< metal1 >>
rect 904 1606 932 1607
rect 904 1603 990 1606
rect 904 1593 908 1603
rect 929 1602 990 1603
rect 929 1601 980 1602
rect 929 1595 934 1601
rect 966 1595 971 1601
rect 904 1592 909 1593
rect 861 1587 909 1592
rect 975 1595 980 1601
rect 885 1580 890 1587
rect 897 1580 902 1587
rect 947 1580 952 1590
rect 947 1576 957 1580
rect 870 1566 875 1575
rect 953 1572 957 1576
rect 916 1569 957 1572
rect 916 1566 919 1569
rect 953 1566 957 1569
rect 859 1562 875 1566
rect 887 1562 919 1566
rect 870 1558 875 1562
rect 927 1561 929 1564
rect 885 1549 890 1553
rect 927 1550 930 1561
rect 944 1558 947 1561
rect 971 1550 974 1564
rect 859 1544 895 1549
rect 859 1543 866 1544
rect 927 1545 974 1550
rect 859 1522 864 1543
rect 936 1535 941 1536
rect 959 1520 964 1536
rect 950 1517 964 1520
rect 809 1510 857 1511
rect 985 1510 990 1602
rect 1247 1510 1270 1511
rect 647 1507 1271 1510
rect 647 1506 1262 1507
rect 647 1505 800 1506
rect 661 1494 666 1505
rect 737 1494 742 1505
rect 759 1498 764 1505
rect 771 1498 776 1505
rect 816 1499 821 1506
rect 828 1499 833 1506
rect 725 1467 730 1489
rect 786 1484 791 1493
rect 843 1485 848 1494
rect 944 1485 948 1493
rect 795 1484 831 1485
rect 756 1480 774 1484
rect 786 1481 831 1484
rect 843 1481 948 1485
rect 786 1480 829 1481
rect 756 1467 759 1480
rect 786 1476 791 1480
rect 843 1477 848 1481
rect 771 1467 776 1471
rect 828 1468 833 1472
rect 819 1467 858 1468
rect 677 1463 759 1467
rect 762 1463 882 1467
rect 677 1458 682 1463
rect 709 1458 714 1463
rect 762 1462 801 1463
rect 889 1463 1181 1467
rect 661 1449 666 1453
rect 693 1450 698 1453
rect 725 1450 730 1453
rect 762 1450 767 1462
rect 693 1449 767 1450
rect 661 1446 767 1449
rect 669 1433 674 1435
rect 685 1431 690 1435
rect 685 1418 689 1431
rect 701 1430 706 1435
rect 722 1436 866 1437
rect 717 1432 866 1436
rect 1178 1436 1181 1463
rect 1266 1454 1271 1507
rect 685 1415 795 1418
rect 292 1406 934 1408
rect 292 1405 935 1406
rect 292 1341 295 1405
rect 655 1382 660 1397
rect 796 1382 800 1397
rect 931 1384 935 1405
rect 141 1338 295 1341
rect 178 1337 295 1338
rect 578 1370 585 1373
rect 928 1370 952 1371
rect 578 1367 1066 1370
rect 94 1315 186 1317
rect 93 1310 186 1315
rect 76 887 82 1296
rect 77 886 82 887
rect 93 1077 99 1310
rect 460 1296 461 1302
rect 475 1296 554 1302
rect 379 1283 530 1288
rect 178 1279 372 1283
rect 178 1245 183 1279
rect 193 1267 356 1271
rect 193 1266 308 1267
rect 193 1259 198 1266
rect 205 1259 210 1266
rect 279 1259 284 1266
rect 220 1245 225 1254
rect 291 1259 296 1266
rect 303 1255 308 1266
rect 178 1242 208 1245
rect 204 1241 208 1242
rect 220 1241 229 1245
rect 264 1245 269 1254
rect 315 1255 320 1267
rect 238 1241 269 1245
rect 281 1241 287 1245
rect 220 1237 225 1241
rect 205 1228 210 1232
rect 196 1223 227 1228
rect 238 1177 242 1241
rect 264 1237 269 1241
rect 294 1241 302 1245
rect 298 1238 302 1241
rect 349 1244 354 1250
rect 367 1244 372 1279
rect 379 1281 384 1283
rect 398 1261 451 1267
rect 398 1255 403 1261
rect 432 1244 437 1250
rect 349 1239 437 1244
rect 298 1233 319 1238
rect 279 1228 284 1232
rect 255 1223 293 1228
rect 283 1186 288 1223
rect 349 1216 354 1239
rect 304 1205 309 1208
rect 383 1215 389 1228
rect 315 1186 320 1211
rect 398 1216 403 1226
rect 432 1216 437 1239
rect 446 1186 451 1261
rect 463 1223 506 1228
rect 465 1216 470 1223
rect 477 1216 482 1223
rect 492 1203 497 1211
rect 511 1203 516 1283
rect 548 1213 554 1296
rect 578 1248 585 1367
rect 717 1357 736 1362
rect 607 1231 611 1356
rect 655 1319 660 1356
rect 717 1321 725 1357
rect 796 1321 800 1359
rect 853 1327 889 1334
rect 717 1320 743 1321
rect 717 1318 744 1320
rect 736 1316 744 1318
rect 690 1310 722 1315
rect 736 1314 738 1316
rect 882 1318 888 1327
rect 883 1317 888 1318
rect 899 1317 904 1322
rect 931 1316 935 1358
rect 1061 1318 1066 1367
rect 1077 1336 1081 1386
rect 1178 1328 1182 1436
rect 1265 1434 1271 1454
rect 1077 1318 1081 1325
rect 617 1303 1130 1307
rect 1265 1305 1270 1434
rect 2097 1359 2104 1360
rect 2097 1355 2362 1359
rect 2097 1354 2370 1355
rect 2071 1335 2076 1340
rect 2097 1335 2104 1354
rect 2071 1329 2104 1335
rect 1248 1304 1349 1305
rect 618 1302 666 1303
rect 642 1295 647 1302
rect 654 1295 659 1302
rect 698 1291 703 1303
rect 730 1291 735 1303
rect 762 1291 767 1303
rect 807 1302 855 1303
rect 627 1281 632 1290
rect 831 1295 836 1302
rect 682 1283 687 1286
rect 714 1283 719 1286
rect 682 1282 719 1283
rect 746 1282 751 1286
rect 622 1277 632 1281
rect 644 1278 668 1281
rect 644 1277 659 1278
rect 627 1273 632 1277
rect 642 1264 647 1268
rect 664 1269 668 1278
rect 682 1278 751 1282
rect 796 1281 800 1291
rect 843 1295 848 1302
rect 863 1291 868 1303
rect 816 1281 821 1290
rect 875 1291 880 1303
rect 907 1291 912 1303
rect 939 1291 944 1303
rect 965 1302 1130 1303
rect 989 1295 994 1302
rect 1001 1295 1006 1302
rect 1027 1290 1032 1302
rect 1053 1290 1058 1302
rect 1085 1290 1090 1302
rect 891 1283 896 1286
rect 876 1282 896 1283
rect 923 1282 928 1286
rect 682 1269 687 1278
rect 796 1277 821 1281
rect 833 1277 852 1281
rect 664 1264 687 1269
rect 816 1273 821 1277
rect 831 1264 836 1268
rect 848 1269 852 1277
rect 876 1278 928 1282
rect 876 1269 881 1278
rect 974 1281 979 1290
rect 1036 1285 1037 1290
rect 1124 1289 1130 1302
rect 1163 1303 1194 1304
rect 1241 1303 1349 1304
rect 1163 1300 1349 1303
rect 1167 1289 1171 1300
rect 1036 1282 1042 1285
rect 1069 1282 1074 1285
rect 1123 1284 1171 1289
rect 1191 1298 1242 1300
rect 1248 1299 1349 1300
rect 1191 1292 1196 1298
rect 1228 1292 1233 1298
rect 1237 1292 1242 1298
rect 967 1277 979 1281
rect 991 1277 1017 1281
rect 1036 1277 1074 1282
rect 1147 1277 1152 1284
rect 848 1264 881 1269
rect 974 1273 979 1277
rect 989 1264 994 1268
rect 1013 1264 1017 1277
rect 1034 1264 1039 1277
rect 1159 1277 1164 1284
rect 1209 1277 1214 1287
rect 1209 1273 1219 1277
rect 617 1259 656 1264
rect 651 1243 656 1259
rect 682 1257 687 1264
rect 806 1259 845 1264
rect 762 1245 767 1252
rect 840 1245 845 1259
rect 876 1257 881 1264
rect 963 1259 1009 1264
rect 1013 1259 1039 1264
rect 762 1243 845 1245
rect 939 1250 944 1252
rect 964 1250 970 1259
rect 939 1247 970 1250
rect 1005 1258 1009 1259
rect 939 1246 949 1247
rect 939 1243 944 1246
rect 651 1240 944 1243
rect 1005 1244 1010 1258
rect 1034 1256 1039 1259
rect 1132 1263 1137 1272
rect 1215 1269 1219 1273
rect 1178 1266 1219 1269
rect 1178 1263 1181 1266
rect 1215 1263 1219 1266
rect 1126 1259 1137 1263
rect 1149 1259 1181 1263
rect 1085 1244 1090 1251
rect 1132 1255 1137 1259
rect 1189 1258 1191 1261
rect 1147 1246 1152 1250
rect 1189 1247 1192 1258
rect 1206 1255 1209 1258
rect 1233 1247 1236 1261
rect 1121 1244 1157 1246
rect 1005 1241 1157 1244
rect 1005 1240 1130 1241
rect 1189 1242 1236 1247
rect 651 1239 767 1240
rect 840 1239 944 1240
rect 607 1229 690 1231
rect 607 1227 695 1229
rect 706 1222 711 1229
rect 754 1226 759 1229
rect 706 1218 737 1222
rect 548 1211 683 1213
rect 548 1208 684 1211
rect 477 1198 480 1202
rect 492 1198 516 1203
rect 492 1194 497 1198
rect 678 1194 684 1208
rect 728 1207 736 1218
rect 730 1199 736 1207
rect 753 1213 762 1226
rect 915 1225 920 1229
rect 1045 1226 1049 1229
rect 753 1206 755 1213
rect 728 1198 736 1199
rect 283 1185 451 1186
rect 477 1185 482 1189
rect 283 1181 530 1185
rect 446 1180 530 1181
rect 238 1172 407 1177
rect 402 1167 407 1172
rect 424 1167 429 1171
rect 402 1162 429 1167
rect 93 1074 224 1077
rect 93 1073 99 1074
rect 93 886 98 1073
rect 507 1066 514 1132
rect 376 1061 514 1066
rect 175 1057 369 1061
rect 175 1023 180 1057
rect 190 1045 353 1049
rect 190 1044 305 1045
rect 190 1037 195 1044
rect 202 1037 207 1044
rect 276 1037 281 1044
rect 217 1023 222 1032
rect 288 1037 293 1044
rect 300 1033 305 1044
rect 175 1020 205 1023
rect 201 1019 205 1020
rect 217 1019 226 1023
rect 261 1023 266 1032
rect 312 1033 317 1045
rect 235 1019 266 1023
rect 278 1021 299 1023
rect 278 1019 286 1021
rect 217 1015 222 1019
rect 202 1006 207 1010
rect 193 1001 224 1006
rect 235 955 239 1019
rect 261 1015 266 1019
rect 292 1019 299 1021
rect 295 1016 299 1019
rect 346 1022 351 1028
rect 364 1022 369 1057
rect 376 1059 381 1061
rect 395 1039 448 1045
rect 395 1033 400 1039
rect 429 1022 434 1028
rect 346 1017 434 1022
rect 295 1011 316 1016
rect 276 1006 281 1010
rect 252 1001 290 1006
rect 280 964 285 1001
rect 346 994 351 1017
rect 395 1011 398 1014
rect 388 1006 403 1011
rect 301 983 306 986
rect 380 995 385 1006
rect 395 994 400 1006
rect 429 994 434 1017
rect 312 964 317 989
rect 443 964 448 1039
rect 460 1001 503 1006
rect 462 994 467 1001
rect 474 994 479 1001
rect 489 981 494 989
rect 508 981 513 1061
rect 474 976 477 980
rect 489 976 513 981
rect 523 998 529 1180
rect 548 1143 557 1181
rect 677 1188 684 1194
rect 570 1129 577 1180
rect 620 1156 621 1163
rect 620 1099 627 1156
rect 552 1091 628 1099
rect 677 1091 683 1188
rect 739 1150 748 1175
rect 914 1171 920 1225
rect 1044 1163 1049 1226
rect 1121 1218 1130 1240
rect 1198 1232 1203 1233
rect 1221 1232 1226 1233
rect 1122 1209 1130 1218
rect 1122 1208 1322 1209
rect 1122 1206 1325 1208
rect 1318 1198 1325 1206
rect 739 1144 1109 1150
rect 789 1112 815 1118
rect 1102 1110 1109 1144
rect 727 1095 958 1099
rect 1319 1094 1323 1198
rect 676 1086 683 1091
rect 585 1065 651 1072
rect 677 1043 683 1086
rect 716 1057 747 1058
rect 794 1057 894 1058
rect 716 1056 942 1057
rect 716 1055 1040 1056
rect 1145 1055 1176 1056
rect 1343 1055 1347 1299
rect 1676 1300 1991 1304
rect 1855 1299 1991 1300
rect 2071 1297 2076 1329
rect 2097 1328 2104 1329
rect 2118 1330 2618 1335
rect 2118 1310 2124 1330
rect 2071 1293 2132 1297
rect 2188 1296 2193 1311
rect 2271 1307 2766 1313
rect 2188 1293 2281 1296
rect 1693 1277 1700 1282
rect 2827 1280 2927 1281
rect 2974 1280 3005 1281
rect 2186 1279 2286 1280
rect 2333 1279 2364 1280
rect 2779 1279 3005 1280
rect 2132 1278 2364 1279
rect 2545 1278 2576 1279
rect 2681 1278 3005 1279
rect 1904 1277 1935 1278
rect 2040 1277 2364 1278
rect 2490 1277 3005 1278
rect 1693 1276 2830 1277
rect 1693 1274 2189 1276
rect 1693 1272 1907 1274
rect 1471 1099 1476 1101
rect 1693 1100 1700 1272
rect 1835 1271 1862 1272
rect 1835 1171 1843 1271
rect 1856 1266 1861 1271
rect 1865 1266 1870 1272
rect 1902 1266 1907 1272
rect 1927 1273 2043 1274
rect 1927 1263 1931 1273
rect 1992 1272 2043 1273
rect 1992 1266 1997 1272
rect 1884 1251 1889 1261
rect 1927 1258 1975 1263
rect 2001 1266 2006 1272
rect 2038 1266 2043 1272
rect 2063 1263 2067 1274
rect 2139 1268 2143 1274
rect 2147 1268 2152 1274
rect 2184 1268 2189 1274
rect 2209 1265 2213 1276
rect 2285 1274 2336 1276
rect 2285 1268 2290 1274
rect 1879 1247 1889 1251
rect 1934 1251 1939 1258
rect 1879 1243 1883 1247
rect 1946 1251 1951 1258
rect 2020 1251 2025 1261
rect 2063 1258 2111 1263
rect 1879 1240 1920 1243
rect 1879 1237 1883 1240
rect 1917 1237 1920 1240
rect 1961 1237 1966 1246
rect 2015 1247 2025 1251
rect 2070 1251 2075 1258
rect 2015 1243 2019 1247
rect 2082 1251 2087 1258
rect 2166 1253 2171 1263
rect 2209 1260 2257 1265
rect 2294 1268 2299 1274
rect 2331 1268 2336 1274
rect 2356 1275 2830 1276
rect 2356 1273 2548 1275
rect 2356 1265 2360 1273
rect 2490 1272 2503 1273
rect 2497 1267 2502 1272
rect 2015 1240 2056 1243
rect 1862 1221 1865 1235
rect 1907 1232 1909 1235
rect 1917 1233 1949 1237
rect 1961 1233 1980 1237
rect 1889 1229 1892 1232
rect 1906 1221 1909 1232
rect 1961 1229 1966 1233
rect 2015 1237 2019 1240
rect 2053 1237 2056 1240
rect 2097 1237 2102 1246
rect 2161 1249 2171 1253
rect 2216 1253 2221 1260
rect 2161 1245 2165 1249
rect 2228 1253 2233 1260
rect 2313 1253 2318 1263
rect 2356 1260 2404 1265
rect 2506 1267 2511 1273
rect 2543 1267 2548 1273
rect 2568 1274 2684 1275
rect 2568 1264 2572 1274
rect 2633 1273 2684 1274
rect 2633 1267 2638 1273
rect 2161 1242 2202 1245
rect 2161 1239 2165 1242
rect 2199 1239 2202 1242
rect 2243 1239 2248 1248
rect 2308 1249 2318 1253
rect 2363 1253 2368 1260
rect 2308 1245 2312 1249
rect 2375 1253 2380 1260
rect 2525 1252 2530 1262
rect 2568 1259 2616 1264
rect 2642 1267 2647 1273
rect 2679 1267 2684 1273
rect 2704 1264 2708 1275
rect 2779 1269 2784 1275
rect 2788 1269 2793 1275
rect 2825 1269 2830 1275
rect 2850 1266 2854 1277
rect 2926 1275 2977 1277
rect 2926 1269 2931 1275
rect 2308 1242 2349 1245
rect 1862 1216 1909 1221
rect 1946 1220 1951 1224
rect 1998 1221 2001 1235
rect 2043 1232 2045 1235
rect 2053 1233 2085 1237
rect 2097 1233 2118 1237
rect 2025 1229 2028 1232
rect 2042 1221 2045 1232
rect 2097 1229 2102 1233
rect 1941 1215 1976 1220
rect 1998 1216 2045 1221
rect 1872 1206 1877 1207
rect 1895 1206 1900 1207
rect 1972 1194 1976 1215
rect 2082 1220 2087 1224
rect 2144 1223 2147 1237
rect 2189 1234 2191 1237
rect 2199 1235 2231 1239
rect 2243 1235 2264 1239
rect 2171 1231 2174 1234
rect 2188 1223 2191 1234
rect 2243 1231 2248 1235
rect 2308 1239 2312 1242
rect 2346 1239 2349 1242
rect 2390 1239 2395 1248
rect 2520 1248 2530 1252
rect 2575 1252 2580 1259
rect 2520 1244 2524 1248
rect 2587 1252 2592 1259
rect 2661 1252 2666 1262
rect 2704 1259 2752 1264
rect 2520 1241 2561 1244
rect 2077 1219 2112 1220
rect 2077 1215 2125 1219
rect 2144 1218 2191 1223
rect 2228 1222 2233 1226
rect 2291 1223 2294 1237
rect 2336 1234 2338 1237
rect 2346 1235 2378 1239
rect 2390 1235 2420 1239
rect 2318 1231 2321 1234
rect 2335 1223 2338 1234
rect 2390 1231 2395 1235
rect 2520 1238 2524 1241
rect 2558 1238 2561 1241
rect 2602 1238 2607 1247
rect 2656 1248 2666 1252
rect 2711 1252 2716 1259
rect 2656 1244 2660 1248
rect 2723 1252 2728 1259
rect 2807 1254 2812 1264
rect 2850 1261 2898 1266
rect 2935 1269 2940 1275
rect 2972 1269 2977 1275
rect 2997 1266 3001 1277
rect 2656 1241 2697 1244
rect 2656 1238 2660 1241
rect 2694 1238 2697 1241
rect 2738 1238 2743 1247
rect 2802 1250 2812 1254
rect 2857 1254 2862 1261
rect 2802 1246 2806 1250
rect 2869 1254 2874 1261
rect 2954 1254 2959 1264
rect 2997 1261 3045 1266
rect 2802 1243 2843 1246
rect 2802 1240 2806 1243
rect 2840 1240 2843 1243
rect 2884 1240 2889 1249
rect 2949 1250 2959 1254
rect 3004 1254 3009 1261
rect 2949 1246 2953 1250
rect 3016 1254 3021 1261
rect 2949 1243 2990 1246
rect 2949 1240 2953 1243
rect 2987 1240 2990 1243
rect 3031 1240 3036 1249
rect 2223 1217 2261 1222
rect 2291 1218 2338 1223
rect 2106 1214 2125 1215
rect 2008 1206 2013 1207
rect 2031 1206 2036 1207
rect 2116 1194 2123 1214
rect 2154 1208 2159 1209
rect 2177 1208 2182 1209
rect 2252 1194 2261 1217
rect 2375 1222 2380 1226
rect 2503 1222 2506 1236
rect 2548 1233 2550 1236
rect 2558 1234 2590 1238
rect 2602 1234 2610 1238
rect 2530 1230 2533 1233
rect 2547 1222 2550 1233
rect 2602 1230 2607 1234
rect 2370 1217 2406 1222
rect 2503 1217 2550 1222
rect 2301 1208 2306 1209
rect 2324 1208 2329 1209
rect 2397 1194 2406 1217
rect 2587 1221 2592 1225
rect 2639 1222 2642 1236
rect 2684 1233 2686 1236
rect 2694 1234 2726 1238
rect 2738 1234 2746 1238
rect 2666 1230 2669 1233
rect 2683 1222 2686 1233
rect 2738 1230 2743 1234
rect 2582 1216 2617 1221
rect 2639 1217 2686 1222
rect 2513 1207 2518 1208
rect 2536 1207 2541 1208
rect 2613 1195 2617 1216
rect 2723 1221 2728 1225
rect 2785 1224 2788 1238
rect 2830 1235 2832 1238
rect 2840 1236 2872 1240
rect 2884 1236 2892 1240
rect 2812 1232 2815 1235
rect 2829 1224 2832 1235
rect 2884 1232 2889 1236
rect 2718 1220 2753 1221
rect 2718 1216 2766 1220
rect 2785 1219 2832 1224
rect 2869 1223 2874 1227
rect 2932 1224 2935 1238
rect 2977 1235 2979 1238
rect 2987 1236 3019 1240
rect 3031 1236 3039 1240
rect 2959 1232 2962 1235
rect 2976 1224 2979 1235
rect 3031 1232 3036 1236
rect 2864 1218 2902 1223
rect 2932 1219 2979 1224
rect 2747 1215 2766 1216
rect 2649 1207 2654 1208
rect 2672 1207 2677 1208
rect 2757 1195 2764 1215
rect 2795 1209 2800 1210
rect 2818 1209 2823 1210
rect 2893 1195 2902 1218
rect 3016 1223 3021 1227
rect 3011 1218 3047 1223
rect 2942 1209 2947 1210
rect 2965 1209 2970 1210
rect 3038 1195 3047 1218
rect 2425 1194 2433 1195
rect 1972 1188 2433 1194
rect 2613 1190 3048 1195
rect 2613 1189 3023 1190
rect 2425 1177 2433 1188
rect 2634 1177 2643 1189
rect 2342 1172 2373 1173
rect 2197 1171 2373 1172
rect 1835 1169 1865 1171
rect 2073 1170 2373 1171
rect 1904 1169 1935 1170
rect 2048 1169 2373 1170
rect 2424 1169 2643 1177
rect 1835 1168 2345 1169
rect 1835 1166 2200 1168
rect 2209 1167 2345 1168
rect 1835 1164 1907 1166
rect 1926 1164 2051 1166
rect 1856 1158 1861 1164
rect 1865 1158 1870 1164
rect 1902 1158 1907 1164
rect 1927 1155 1931 1164
rect 2000 1158 2005 1164
rect 1884 1143 1889 1153
rect 1927 1150 1975 1155
rect 2009 1158 2014 1164
rect 2046 1158 2051 1164
rect 2071 1155 2075 1166
rect 2149 1160 2154 1166
rect 2158 1160 2163 1166
rect 2195 1160 2200 1166
rect 2220 1157 2224 1167
rect 2294 1161 2299 1167
rect 1879 1139 1889 1143
rect 1934 1143 1939 1150
rect 1879 1135 1883 1139
rect 1946 1143 1951 1150
rect 2028 1143 2033 1153
rect 2071 1150 2119 1155
rect 1879 1132 1920 1135
rect 1879 1129 1883 1132
rect 1917 1129 1920 1132
rect 1961 1129 1966 1138
rect 2023 1139 2033 1143
rect 2078 1143 2083 1150
rect 2023 1135 2027 1139
rect 2090 1143 2095 1150
rect 2177 1145 2182 1155
rect 2220 1152 2268 1157
rect 2303 1161 2308 1167
rect 2340 1161 2345 1167
rect 2365 1158 2369 1169
rect 2023 1132 2064 1135
rect 1862 1113 1865 1127
rect 1907 1124 1909 1127
rect 1917 1125 1949 1129
rect 1961 1125 1993 1129
rect 1889 1121 1892 1124
rect 1906 1113 1909 1124
rect 1961 1121 1966 1125
rect 2023 1129 2027 1132
rect 2061 1129 2064 1132
rect 2105 1129 2110 1138
rect 2172 1141 2182 1145
rect 2227 1145 2232 1152
rect 2172 1137 2176 1141
rect 2239 1145 2244 1152
rect 2322 1146 2327 1156
rect 2365 1153 2413 1158
rect 2172 1134 2213 1137
rect 2172 1131 2176 1134
rect 2210 1131 2213 1134
rect 2254 1131 2259 1140
rect 2317 1142 2327 1146
rect 2372 1146 2377 1153
rect 2317 1138 2321 1142
rect 2384 1146 2389 1153
rect 2317 1135 2358 1138
rect 2317 1132 2321 1135
rect 2355 1132 2358 1135
rect 2399 1132 2404 1141
rect 1862 1108 1909 1113
rect 1946 1112 1951 1116
rect 2006 1113 2009 1127
rect 2051 1124 2053 1127
rect 2061 1125 2093 1129
rect 2105 1125 2133 1129
rect 2033 1121 2036 1124
rect 2050 1113 2053 1124
rect 2105 1121 2110 1125
rect 1941 1107 1976 1112
rect 2006 1108 2053 1113
rect 1597 1099 1700 1100
rect 1471 1096 1701 1099
rect 1471 1095 1600 1096
rect 1471 1055 1476 1095
rect 1549 1094 1600 1095
rect 1549 1088 1554 1094
rect 1558 1088 1563 1094
rect 1595 1088 1600 1094
rect 1620 1086 1624 1096
rect 1693 1086 1701 1096
rect 1872 1098 1877 1099
rect 1895 1098 1900 1099
rect 1577 1073 1582 1083
rect 1618 1081 1701 1086
rect 1572 1069 1582 1073
rect 1625 1074 1630 1081
rect 1637 1074 1642 1081
rect 1572 1065 1576 1069
rect 1572 1062 1613 1065
rect 1572 1059 1576 1062
rect 1610 1059 1613 1062
rect 1652 1060 1657 1069
rect 1693 1061 1701 1081
rect 1617 1059 1640 1060
rect 716 1054 1476 1055
rect 720 1043 724 1054
rect 676 1038 724 1043
rect 744 1052 795 1054
rect 744 1046 749 1052
rect 781 1046 786 1052
rect 790 1046 795 1052
rect 867 1043 871 1054
rect 700 1031 705 1038
rect 712 1031 717 1038
rect 762 1031 767 1041
rect 823 1038 871 1043
rect 891 1052 1476 1054
rect 891 1046 896 1052
rect 928 1046 933 1052
rect 937 1046 942 1052
rect 1013 1041 1017 1052
rect 847 1031 852 1038
rect 762 1027 772 1031
rect 685 1017 690 1026
rect 768 1023 772 1027
rect 731 1020 772 1023
rect 731 1017 734 1020
rect 768 1017 772 1020
rect 859 1031 864 1038
rect 909 1031 914 1041
rect 969 1036 1017 1041
rect 1037 1051 1153 1052
rect 1037 1050 1088 1051
rect 1037 1044 1042 1050
rect 1074 1044 1079 1050
rect 1083 1044 1088 1050
rect 1149 1041 1153 1051
rect 909 1027 919 1031
rect 993 1029 998 1036
rect 667 1013 690 1017
rect 702 1013 734 1017
rect 685 1009 690 1013
rect 742 1012 744 1015
rect 700 1000 705 1004
rect 742 1001 745 1012
rect 759 1009 762 1012
rect 786 1001 789 1015
rect 832 1017 837 1026
rect 915 1023 919 1027
rect 878 1020 919 1023
rect 878 1017 881 1020
rect 915 1017 919 1020
rect 1005 1029 1010 1036
rect 1055 1029 1060 1039
rect 1105 1036 1153 1041
rect 1173 1050 1476 1052
rect 1173 1044 1178 1050
rect 1210 1044 1215 1050
rect 1218 1049 1476 1050
rect 1219 1044 1224 1049
rect 1129 1029 1134 1036
rect 1055 1025 1065 1029
rect 821 1014 837 1017
rect 819 1013 837 1014
rect 849 1013 881 1017
rect 832 1009 837 1013
rect 889 1012 891 1015
rect 674 998 710 1000
rect 523 995 710 998
rect 523 993 683 995
rect 742 996 789 1001
rect 847 1000 852 1004
rect 889 1001 892 1012
rect 906 1009 909 1012
rect 933 1001 936 1015
rect 978 1015 983 1024
rect 1061 1021 1065 1025
rect 1024 1018 1065 1021
rect 1024 1015 1027 1018
rect 1061 1015 1065 1018
rect 1141 1029 1146 1036
rect 1191 1029 1196 1039
rect 1191 1025 1201 1029
rect 1114 1015 1119 1024
rect 1197 1021 1201 1025
rect 1160 1018 1201 1021
rect 1160 1015 1163 1018
rect 1197 1015 1201 1018
rect 966 1011 983 1015
rect 995 1011 1027 1015
rect 978 1007 983 1011
rect 1035 1010 1037 1013
rect 1104 1014 1119 1015
rect 819 995 857 1000
rect 489 972 494 976
rect 280 963 448 964
rect 474 963 479 967
rect 523 963 529 993
rect 280 959 529 963
rect 443 958 529 959
rect 235 950 404 955
rect 399 945 404 950
rect 421 945 426 949
rect 160 934 198 938
rect 399 940 426 945
rect 160 933 202 934
rect 483 881 488 893
rect 144 876 149 881
rect 379 876 516 881
rect 1 872 149 876
rect 153 872 372 876
rect 1 871 49 872
rect 25 864 30 871
rect 37 864 42 871
rect 57 860 62 872
rect 10 850 15 859
rect 69 860 74 872
rect 101 860 106 872
rect 133 860 138 872
rect 85 852 90 855
rect 70 851 90 852
rect 117 851 122 855
rect 3 846 15 850
rect 27 846 46 850
rect 10 842 15 846
rect 25 833 30 837
rect 42 838 46 846
rect 70 847 122 851
rect 70 838 75 847
rect 42 833 45 838
rect 50 833 75 838
rect 153 838 158 872
rect 168 860 356 864
rect 168 859 308 860
rect 168 852 173 859
rect 205 852 210 859
rect 279 852 284 859
rect 220 838 225 847
rect 291 852 296 859
rect 303 848 308 859
rect 264 838 269 847
rect 315 848 320 860
rect 153 835 208 838
rect 204 834 208 835
rect 220 834 228 838
rect 0 828 39 833
rect 34 812 39 828
rect 70 826 75 833
rect 220 830 225 834
rect 238 834 269 838
rect 281 836 302 838
rect 281 834 288 836
rect 205 821 210 825
rect 133 819 138 821
rect 171 819 227 821
rect 133 816 227 819
rect 133 815 175 816
rect 133 812 138 815
rect 34 808 138 812
rect 153 801 186 804
rect 109 782 114 798
rect 125 793 130 798
rect 125 789 226 793
rect 109 778 143 782
rect 238 770 242 834
rect 264 830 269 834
rect 293 834 302 836
rect 298 831 302 834
rect 349 837 354 843
rect 367 837 372 872
rect 379 874 384 876
rect 398 854 451 860
rect 398 848 403 854
rect 432 837 437 843
rect 349 832 437 837
rect 298 826 319 831
rect 279 821 284 825
rect 255 816 293 821
rect 283 779 288 816
rect 349 809 354 832
rect 398 826 401 829
rect 304 798 309 801
rect 391 821 406 826
rect 383 808 388 821
rect 315 779 320 804
rect 398 809 403 821
rect 432 809 437 832
rect 446 779 451 854
rect 463 816 506 821
rect 465 809 470 816
rect 477 809 482 816
rect 492 796 497 804
rect 511 796 516 876
rect 477 791 480 795
rect 492 791 516 796
rect 492 787 497 791
rect 283 778 451 779
rect 477 778 482 782
rect 523 778 529 958
rect 541 965 542 974
rect 647 972 655 973
rect 674 972 683 993
rect 751 986 756 987
rect 774 986 779 987
rect 819 972 828 995
rect 889 996 936 1001
rect 993 998 998 1002
rect 1035 999 1038 1010
rect 1052 1007 1055 1010
rect 1079 999 1082 1013
rect 1109 1011 1119 1014
rect 1131 1011 1163 1015
rect 1114 1007 1119 1011
rect 1171 1010 1173 1013
rect 968 997 1003 998
rect 955 993 1003 997
rect 898 986 903 987
rect 955 992 974 993
rect 1035 994 1082 999
rect 1129 998 1134 1002
rect 1171 999 1174 1010
rect 1188 1007 1191 1010
rect 1215 999 1218 1013
rect 1104 993 1139 998
rect 921 986 926 987
rect 957 972 964 992
rect 1044 984 1049 985
rect 1067 984 1072 985
rect 1104 972 1108 993
rect 1171 994 1218 999
rect 1180 984 1185 985
rect 1203 984 1208 985
rect 541 922 548 965
rect 575 888 581 971
rect 647 966 1108 972
rect 545 882 581 888
rect 618 857 620 866
rect 618 789 627 857
rect 283 774 531 778
rect 446 773 531 774
rect 238 765 407 770
rect 402 760 407 765
rect 424 760 429 764
rect 402 755 429 760
rect 502 736 506 758
rect 379 701 510 706
rect 178 697 372 701
rect 178 663 183 697
rect 193 685 356 689
rect 193 684 308 685
rect 193 677 198 684
rect 205 677 210 684
rect 279 677 284 684
rect 220 663 225 672
rect 291 677 296 684
rect 303 673 308 684
rect 264 663 269 672
rect 315 673 320 685
rect 178 660 208 663
rect 204 659 208 660
rect 220 659 228 663
rect 220 655 225 659
rect 238 659 269 663
rect 281 661 302 663
rect 281 659 288 661
rect 205 646 210 650
rect 196 641 227 646
rect 238 595 242 659
rect 264 655 269 659
rect 294 659 302 661
rect 298 656 302 659
rect 349 662 354 668
rect 367 662 372 697
rect 379 699 384 701
rect 398 679 451 685
rect 398 673 403 679
rect 432 662 437 668
rect 349 657 437 662
rect 298 651 319 656
rect 279 646 284 650
rect 255 641 293 646
rect 283 604 288 641
rect 349 634 354 657
rect 398 651 401 654
rect 388 646 406 651
rect 304 623 309 626
rect 379 634 386 646
rect 398 634 403 646
rect 379 629 383 634
rect 432 634 437 657
rect 315 604 320 629
rect 446 604 451 679
rect 463 641 506 646
rect 465 634 470 641
rect 477 634 482 641
rect 492 621 497 629
rect 511 621 516 701
rect 477 616 480 620
rect 492 616 516 621
rect 492 612 497 616
rect 283 603 451 604
rect 477 603 482 607
rect 523 603 529 773
rect 617 705 627 789
rect 617 640 626 705
rect 283 599 529 603
rect 446 598 529 599
rect 238 590 407 595
rect 402 585 407 590
rect 424 585 429 589
rect 402 580 429 585
rect 476 562 483 571
rect 635 562 641 906
rect 647 860 655 966
rect 707 950 738 951
rect 707 949 883 950
rect 1237 949 1245 1049
rect 707 948 1007 949
rect 707 947 1032 948
rect 1145 947 1176 948
rect 1215 947 1245 949
rect 1471 947 1476 1049
rect 1555 1043 1558 1057
rect 1600 1054 1602 1057
rect 1610 1056 1640 1059
rect 1652 1056 1660 1060
rect 1610 1055 1637 1056
rect 1582 1051 1585 1054
rect 1599 1043 1602 1054
rect 1652 1052 1657 1056
rect 1694 1056 1700 1061
rect 1834 1056 1837 1086
rect 1968 1083 1977 1107
rect 2090 1112 2095 1116
rect 2155 1115 2158 1129
rect 2200 1126 2202 1129
rect 2210 1127 2242 1131
rect 2254 1127 2282 1131
rect 2182 1123 2185 1126
rect 2199 1115 2202 1126
rect 2254 1123 2259 1127
rect 2085 1107 2126 1112
rect 2155 1110 2202 1115
rect 2239 1114 2244 1118
rect 2300 1116 2303 1130
rect 2345 1127 2347 1130
rect 2355 1128 2387 1132
rect 2399 1128 2407 1132
rect 2327 1124 2330 1127
rect 2344 1116 2347 1127
rect 2399 1124 2404 1128
rect 2234 1109 2269 1114
rect 2300 1111 2347 1116
rect 2384 1115 2389 1119
rect 2408 1115 2415 1116
rect 2379 1110 2415 1115
rect 2016 1098 2021 1099
rect 2039 1098 2044 1099
rect 2118 1083 2125 1107
rect 2165 1100 2170 1101
rect 2188 1100 2193 1101
rect 2262 1083 2269 1109
rect 2310 1100 2315 1102
rect 2333 1101 2338 1102
rect 2408 1083 2415 1110
rect 1968 1082 2415 1083
rect 2425 1082 2433 1169
rect 2634 1168 2643 1169
rect 1968 1077 2433 1082
rect 1637 1043 1642 1047
rect 1555 1038 1602 1043
rect 1634 1038 1656 1043
rect 1649 1037 1656 1038
rect 711 936 715 947
rect 667 931 715 936
rect 735 946 1245 947
rect 735 945 871 946
rect 735 939 740 945
rect 772 939 777 945
rect 781 939 786 945
rect 856 935 860 945
rect 691 924 696 931
rect 703 924 708 931
rect 753 924 758 934
rect 812 930 860 935
rect 880 944 1245 946
rect 880 938 885 944
rect 917 938 922 944
rect 926 938 931 944
rect 1005 933 1009 944
rect 753 920 763 924
rect 836 923 841 930
rect 676 910 681 919
rect 759 916 763 920
rect 722 913 763 916
rect 722 910 725 913
rect 759 910 763 913
rect 848 923 853 930
rect 898 923 903 933
rect 961 928 1009 933
rect 1029 942 1154 944
rect 1173 942 1245 944
rect 1390 942 1476 947
rect 1693 1042 1701 1056
rect 1692 1037 1702 1042
rect 1029 936 1034 942
rect 1066 936 1071 942
rect 1075 936 1080 942
rect 1149 933 1153 942
rect 898 919 908 923
rect 985 921 990 928
rect 668 906 681 910
rect 693 906 725 910
rect 676 902 681 906
rect 733 905 735 908
rect 665 893 672 894
rect 691 893 696 897
rect 733 894 736 905
rect 750 902 753 905
rect 777 894 780 908
rect 821 909 826 918
rect 904 915 908 919
rect 867 912 908 915
rect 867 909 870 912
rect 904 909 908 912
rect 997 921 1002 928
rect 1047 921 1052 931
rect 1105 928 1153 933
rect 1173 936 1178 942
rect 1210 936 1215 942
rect 1219 936 1224 942
rect 1397 935 1402 942
rect 1129 921 1134 928
rect 1047 917 1057 921
rect 809 906 826 909
rect 818 905 826 906
rect 838 905 870 909
rect 821 901 826 905
rect 878 904 880 907
rect 970 907 975 916
rect 1053 913 1057 917
rect 1016 910 1057 913
rect 1016 907 1019 910
rect 1053 907 1057 910
rect 1141 921 1146 928
rect 1191 921 1196 931
rect 1409 935 1414 942
rect 1447 935 1452 942
rect 1191 917 1201 921
rect 665 888 701 893
rect 665 861 672 888
rect 733 889 780 894
rect 836 892 841 896
rect 878 893 881 904
rect 895 901 898 904
rect 922 893 925 907
rect 952 902 975 907
rect 987 903 1019 907
rect 970 899 975 902
rect 1027 902 1029 905
rect 811 887 846 892
rect 742 879 747 880
rect 765 878 770 880
rect 811 861 818 887
rect 878 888 925 893
rect 985 890 990 894
rect 1027 891 1030 902
rect 1044 899 1047 902
rect 1071 891 1074 905
rect 1114 907 1119 916
rect 1197 913 1201 917
rect 1410 917 1412 921
rect 1410 916 1411 917
rect 1424 913 1429 930
rect 1462 921 1467 930
rect 1447 917 1450 921
rect 1462 916 1465 921
rect 1462 913 1467 916
rect 1160 910 1201 913
rect 1160 907 1163 910
rect 1197 907 1201 910
rect 1095 903 1119 907
rect 1131 903 1163 907
rect 1114 899 1119 903
rect 1171 902 1173 905
rect 954 885 995 890
rect 887 878 892 879
rect 910 878 915 879
rect 955 861 962 885
rect 1027 886 1074 891
rect 1129 890 1134 894
rect 1171 891 1174 902
rect 1188 899 1191 902
rect 1215 891 1218 905
rect 1409 904 1414 908
rect 1447 906 1452 908
rect 1434 904 1453 906
rect 1353 903 1479 904
rect 1353 899 1437 903
rect 1450 901 1479 903
rect 1452 899 1479 901
rect 1353 896 1404 899
rect 1104 885 1139 890
rect 1036 876 1041 877
rect 1059 876 1064 877
rect 1103 861 1112 885
rect 1171 886 1218 891
rect 1180 876 1185 877
rect 1203 876 1208 877
rect 1249 868 1318 872
rect 665 860 1112 861
rect 647 855 1112 860
rect 665 854 672 855
rect 955 853 962 855
rect 1103 836 1111 855
rect 1398 836 1404 896
rect 1103 832 1405 836
rect 1319 664 1323 704
rect 1398 694 1404 832
rect 1442 795 1446 894
rect 1488 807 1496 1015
rect 1596 981 1627 982
rect 1548 978 1627 981
rect 1548 976 1599 978
rect 1548 970 1553 976
rect 1557 970 1562 976
rect 1594 970 1599 976
rect 1619 967 1623 978
rect 1693 967 1701 1037
rect 1935 1042 1944 1044
rect 1729 1037 1944 1042
rect 1576 955 1581 965
rect 1617 962 1701 967
rect 1571 951 1581 955
rect 1624 955 1629 962
rect 1571 947 1575 951
rect 1636 955 1641 962
rect 1674 961 1688 962
rect 1571 944 1612 947
rect 1571 941 1575 944
rect 1609 941 1612 944
rect 1651 941 1656 950
rect 1554 925 1557 939
rect 1599 936 1601 939
rect 1609 937 1639 941
rect 1651 937 1666 941
rect 1581 933 1584 936
rect 1598 925 1601 936
rect 1651 933 1656 937
rect 1554 920 1601 925
rect 1636 924 1641 928
rect 1632 919 1662 924
rect 1564 908 1569 911
rect 1586 908 1592 911
rect 1693 913 1701 962
rect 1792 960 1796 1018
rect 1855 1009 1891 1014
rect 1888 993 1891 1009
rect 1935 1008 1944 1037
rect 2076 1008 2083 1077
rect 2118 1075 2125 1077
rect 2408 1076 2415 1077
rect 1935 1002 2084 1008
rect 2076 1000 2083 1002
rect 2162 998 2388 1000
rect 2162 997 2383 998
rect 2162 993 2165 997
rect 1888 990 2165 993
rect 2587 991 2687 992
rect 2734 991 2765 992
rect 2539 990 2765 991
rect 2305 989 2336 990
rect 2441 989 2765 990
rect 2236 988 2765 989
rect 2236 986 2590 988
rect 2236 984 2308 986
rect 2236 983 2263 984
rect 1792 957 2222 960
rect 1738 941 2032 942
rect 1738 940 2042 941
rect 1738 937 2036 940
rect 2024 934 2036 937
rect 2218 932 2222 957
rect 2236 914 2244 983
rect 2257 978 2262 983
rect 2266 978 2271 984
rect 2303 978 2308 984
rect 2328 985 2444 986
rect 2328 975 2332 985
rect 2393 984 2444 985
rect 2393 978 2398 984
rect 2285 963 2290 973
rect 2328 970 2376 975
rect 2402 978 2407 984
rect 2439 978 2444 984
rect 2464 975 2468 986
rect 2539 980 2544 986
rect 2548 980 2553 986
rect 2585 980 2590 986
rect 2610 977 2614 988
rect 2686 986 2737 988
rect 2686 980 2691 986
rect 2280 959 2290 963
rect 2335 963 2340 970
rect 2280 955 2284 959
rect 2347 963 2352 970
rect 2421 963 2426 973
rect 2464 970 2512 975
rect 2280 952 2321 955
rect 2280 949 2284 952
rect 2318 949 2321 952
rect 2362 949 2367 958
rect 2416 959 2426 963
rect 2471 963 2476 970
rect 2416 955 2420 959
rect 2483 963 2488 970
rect 2567 965 2572 975
rect 2610 972 2658 977
rect 2695 980 2700 986
rect 2732 980 2737 986
rect 2757 977 2761 988
rect 2416 952 2457 955
rect 2263 933 2266 947
rect 2308 944 2310 947
rect 2318 945 2350 949
rect 2362 947 2373 949
rect 2416 949 2420 952
rect 2454 949 2457 952
rect 2498 949 2503 958
rect 2562 961 2572 965
rect 2617 965 2622 972
rect 2562 957 2566 961
rect 2629 965 2634 972
rect 2714 965 2719 975
rect 2757 972 2805 977
rect 2562 954 2603 957
rect 2562 951 2566 954
rect 2600 951 2603 954
rect 2644 952 2649 960
rect 2709 961 2719 965
rect 2764 965 2769 972
rect 2709 957 2713 961
rect 2776 965 2781 972
rect 2709 954 2750 957
rect 2362 945 2377 947
rect 2290 941 2293 944
rect 2307 933 2310 944
rect 2362 941 2367 945
rect 2263 928 2310 933
rect 2347 932 2352 936
rect 2399 933 2402 947
rect 2444 944 2446 947
rect 2454 945 2486 949
rect 2498 945 2506 949
rect 2426 941 2429 944
rect 2443 933 2446 944
rect 2498 941 2503 945
rect 2342 927 2377 932
rect 2399 928 2446 933
rect 2055 913 2244 914
rect 1693 909 2244 913
rect 2273 918 2278 919
rect 2296 918 2301 919
rect 1693 908 2055 909
rect 1595 877 1626 878
rect 1547 874 1626 877
rect 1547 872 1598 874
rect 1547 866 1552 872
rect 1556 866 1561 872
rect 1593 866 1598 872
rect 1618 863 1622 874
rect 1693 863 1701 908
rect 1995 900 2000 908
rect 1769 895 1984 899
rect 2005 900 2010 908
rect 2062 902 2067 909
rect 2024 895 2029 900
rect 2074 902 2079 909
rect 1980 885 1984 895
rect 1980 881 2008 885
rect 2004 880 2008 881
rect 2043 884 2048 895
rect 2089 888 2094 897
rect 2061 884 2077 888
rect 2089 884 2099 888
rect 2043 879 2065 884
rect 2089 880 2094 884
rect 2043 877 2048 879
rect 1575 851 1580 861
rect 1618 858 1701 863
rect 2005 871 2048 877
rect 2236 883 2244 909
rect 2373 906 2377 927
rect 2483 932 2488 936
rect 2545 935 2548 949
rect 2590 946 2592 949
rect 2600 947 2632 951
rect 2644 947 2648 952
rect 2709 951 2713 954
rect 2747 951 2750 954
rect 2791 951 2796 960
rect 2572 943 2575 946
rect 2589 935 2592 946
rect 2644 943 2649 947
rect 2478 931 2513 932
rect 2478 927 2526 931
rect 2545 930 2592 935
rect 2629 934 2634 938
rect 2692 935 2695 949
rect 2737 946 2739 949
rect 2747 947 2779 951
rect 2791 947 2818 951
rect 2719 943 2722 946
rect 2736 935 2739 946
rect 2791 943 2796 947
rect 2624 929 2662 934
rect 2692 930 2739 935
rect 2507 926 2526 927
rect 2409 918 2414 919
rect 2432 918 2437 919
rect 2517 906 2524 926
rect 2555 920 2560 921
rect 2578 920 2583 921
rect 2653 906 2662 929
rect 2776 934 2781 938
rect 2771 929 2807 934
rect 2702 920 2707 921
rect 2725 920 2730 921
rect 2798 906 2807 929
rect 2826 906 2834 907
rect 2373 900 2834 906
rect 2743 884 2774 885
rect 2598 883 2774 884
rect 2236 881 2266 883
rect 2474 882 2774 883
rect 2305 881 2336 882
rect 2449 881 2774 882
rect 2236 880 2746 881
rect 2236 878 2601 880
rect 2610 879 2746 880
rect 2236 876 2308 878
rect 2327 876 2452 878
rect 2074 871 2079 875
rect 2005 863 2010 871
rect 2043 863 2048 871
rect 2065 870 2104 871
rect 2257 870 2262 876
rect 2065 866 2243 870
rect 1570 847 1580 851
rect 1625 851 1630 858
rect 1570 843 1574 847
rect 1637 851 1642 858
rect 1570 840 1611 843
rect 1570 837 1574 840
rect 1608 837 1611 840
rect 1652 837 1657 846
rect 1553 821 1556 835
rect 1598 832 1600 835
rect 1608 833 1640 837
rect 1652 833 1670 837
rect 1580 829 1583 832
rect 1597 821 1600 832
rect 1652 829 1657 833
rect 1553 816 1600 821
rect 1637 820 1642 824
rect 1631 815 1658 820
rect 1488 802 1568 807
rect 1586 795 1591 807
rect 1442 789 1591 795
rect 1533 712 1537 789
rect 1595 781 1626 782
rect 1555 778 1626 781
rect 1555 776 1598 778
rect 1547 770 1552 776
rect 1556 770 1561 776
rect 1593 770 1598 776
rect 1618 767 1622 778
rect 1693 767 1701 858
rect 2023 852 2028 858
rect 2065 852 2070 866
rect 2100 865 2243 866
rect 2266 870 2271 876
rect 2303 870 2308 876
rect 2328 867 2332 876
rect 2401 870 2406 876
rect 2023 849 2070 852
rect 2028 845 2032 849
rect 1616 766 1701 767
rect 2019 842 2032 845
rect 1575 755 1580 765
rect 1616 762 2002 766
rect 1570 751 1580 755
rect 1624 755 1629 762
rect 1570 747 1574 751
rect 1636 755 1641 762
rect 1687 761 2002 762
rect 1570 744 1611 747
rect 1570 741 1574 744
rect 1608 741 1611 744
rect 1651 741 1656 750
rect 1553 725 1556 739
rect 1598 736 1600 739
rect 1608 737 1639 741
rect 1651 737 1805 741
rect 1580 733 1583 736
rect 1597 725 1600 736
rect 1651 733 1656 737
rect 1553 720 1600 725
rect 1636 724 1641 728
rect 1657 724 1665 725
rect 1632 719 1665 724
rect 1657 718 1665 719
rect 1774 718 1938 721
rect 1533 711 1563 712
rect 1533 708 1568 711
rect 1659 694 1665 718
rect 1398 693 1665 694
rect 1398 689 2006 693
rect 2019 693 2023 842
rect 2238 787 2243 865
rect 2285 855 2290 865
rect 2328 862 2376 867
rect 2410 870 2415 876
rect 2447 870 2452 876
rect 2472 867 2476 878
rect 2550 872 2555 878
rect 2559 872 2564 878
rect 2596 872 2601 878
rect 2621 869 2625 879
rect 2695 873 2700 879
rect 2280 851 2290 855
rect 2335 855 2340 862
rect 2280 847 2284 851
rect 2347 855 2352 862
rect 2429 855 2434 865
rect 2472 862 2520 867
rect 2280 844 2321 847
rect 2280 841 2284 844
rect 2318 841 2321 844
rect 2263 825 2266 839
rect 2308 836 2310 839
rect 2318 837 2350 841
rect 2290 833 2293 836
rect 2307 825 2310 836
rect 2362 833 2367 850
rect 2424 851 2434 855
rect 2479 855 2484 862
rect 2424 847 2428 851
rect 2491 855 2496 862
rect 2578 857 2583 867
rect 2621 864 2669 869
rect 2704 873 2709 879
rect 2741 873 2746 879
rect 2766 870 2770 881
rect 2424 844 2465 847
rect 2424 841 2428 844
rect 2462 841 2465 844
rect 2506 841 2511 850
rect 2573 853 2583 857
rect 2628 857 2633 864
rect 2573 849 2577 853
rect 2640 857 2645 864
rect 2723 858 2728 868
rect 2766 865 2814 870
rect 2573 846 2614 849
rect 2573 843 2577 846
rect 2611 843 2614 846
rect 2655 843 2660 852
rect 2718 854 2728 858
rect 2773 858 2778 865
rect 2718 850 2722 854
rect 2785 858 2790 865
rect 2718 847 2759 850
rect 2718 844 2722 847
rect 2756 844 2759 847
rect 2800 844 2805 853
rect 2263 820 2310 825
rect 2347 824 2352 828
rect 2407 825 2410 839
rect 2452 836 2454 839
rect 2462 837 2494 841
rect 2506 837 2520 841
rect 2434 833 2437 836
rect 2451 825 2454 836
rect 2506 833 2511 837
rect 2342 819 2377 824
rect 2407 820 2454 825
rect 2273 810 2278 811
rect 2296 810 2301 811
rect 2369 795 2378 819
rect 2491 824 2496 828
rect 2556 827 2559 841
rect 2601 838 2603 841
rect 2611 839 2643 843
rect 2655 839 2667 843
rect 2583 835 2586 838
rect 2600 827 2603 838
rect 2655 835 2660 839
rect 2486 819 2527 824
rect 2556 822 2603 827
rect 2640 826 2645 830
rect 2701 828 2704 842
rect 2746 839 2748 842
rect 2756 840 2788 844
rect 2800 840 2812 844
rect 2728 836 2731 839
rect 2745 828 2748 839
rect 2800 836 2805 840
rect 2635 821 2670 826
rect 2701 823 2748 828
rect 2785 827 2790 831
rect 2809 827 2816 828
rect 2780 822 2816 827
rect 2417 810 2422 811
rect 2440 810 2445 811
rect 2519 795 2526 819
rect 2566 812 2571 813
rect 2589 812 2594 813
rect 2663 795 2670 821
rect 2711 812 2716 814
rect 2734 813 2739 814
rect 2809 795 2816 822
rect 2369 794 2816 795
rect 2826 794 2834 900
rect 2369 789 2834 794
rect 2369 787 2375 789
rect 2519 787 2526 789
rect 2809 788 2816 789
rect 2238 784 2375 787
rect 2011 689 2023 693
rect 2135 671 2272 676
rect 2135 669 2140 671
rect 1319 659 1831 664
rect 2007 655 2036 659
rect 2042 655 2112 659
rect 2007 654 2055 655
rect 2031 647 2036 654
rect 2043 647 2048 654
rect 2059 643 2064 655
rect 2016 633 2021 642
rect 2071 643 2076 655
rect 2154 649 2207 655
rect 2154 643 2159 649
rect 1994 629 2021 633
rect 2033 629 2046 633
rect 476 556 641 562
rect 673 539 682 625
rect 1994 565 1998 629
rect 2016 625 2021 629
rect 2051 629 2058 633
rect 2054 626 2058 629
rect 2105 632 2110 638
rect 2105 627 2122 632
rect 2188 632 2193 638
rect 2128 627 2193 632
rect 2054 621 2075 626
rect 2031 616 2036 620
rect 2012 611 2045 616
rect 2039 574 2044 611
rect 2105 604 2110 627
rect 2154 621 2157 624
rect 2145 616 2162 621
rect 2060 593 2065 596
rect 2139 602 2144 616
rect 2071 574 2076 599
rect 2154 604 2159 616
rect 2188 604 2193 627
rect 2202 574 2207 649
rect 2219 611 2262 616
rect 2221 604 2226 611
rect 2233 604 2238 611
rect 2248 591 2253 599
rect 2267 591 2272 671
rect 2233 586 2236 590
rect 2248 586 2272 591
rect 2248 582 2253 586
rect 2039 573 2207 574
rect 2233 573 2238 577
rect 2039 569 2263 573
rect 2202 568 2263 569
rect 1994 560 2163 565
rect 2158 555 2163 560
rect 2180 555 2185 559
rect 1465 551 1601 553
rect 1465 548 2028 551
rect 2158 550 2185 555
rect 1483 541 1488 548
rect 299 533 682 539
rect 1495 541 1500 548
rect 1522 537 1527 548
rect 1579 537 1584 548
rect 1468 527 1473 536
rect 1595 545 2028 548
rect 1422 523 1473 527
rect 1485 523 1511 527
rect 1468 519 1473 523
rect 1156 510 1163 512
rect 1213 510 1472 511
rect 1483 510 1488 514
rect 1508 510 1511 523
rect 1531 510 1536 532
rect 1156 506 1505 510
rect 1508 506 1568 510
rect 1156 505 1229 506
rect 1458 505 1505 506
rect 1156 -10 1163 505
rect 1500 493 1505 505
rect 1531 501 1536 506
rect 1563 501 1568 506
rect 1547 493 1552 496
rect 1500 492 1552 493
rect 1579 493 1584 496
rect 1500 489 1579 492
rect 1539 477 1544 478
rect 1555 476 1560 478
rect 1571 476 1576 478
rect 1328 434 1356 435
rect 1328 433 1404 434
rect 1328 432 1502 433
rect 1595 432 1601 545
rect 2023 476 2027 545
rect 2129 488 2266 493
rect 2129 486 2134 488
rect 2001 472 2106 476
rect 2001 471 2049 472
rect 2025 464 2030 471
rect 2053 460 2058 472
rect 2010 450 2015 459
rect 2065 460 2070 472
rect 2148 466 2201 472
rect 2148 460 2153 466
rect 1988 446 2015 450
rect 2027 446 2038 450
rect 2043 446 2052 450
rect 1831 436 1841 444
rect 1607 432 1638 433
rect 1832 432 1841 436
rect 1328 431 1841 432
rect 1329 420 1333 431
rect 1259 416 1333 420
rect 1353 429 1841 431
rect 1353 423 1358 429
rect 1390 423 1395 429
rect 1399 423 1404 429
rect 1475 418 1479 429
rect 1184 379 1239 385
rect 1184 6 1188 379
rect 1234 331 1239 379
rect 1259 316 1265 416
rect 1285 415 1333 416
rect 1309 408 1314 415
rect 1321 408 1326 415
rect 1371 408 1376 418
rect 1431 413 1479 418
rect 1499 428 1615 429
rect 1499 427 1550 428
rect 1499 421 1504 427
rect 1536 421 1541 427
rect 1545 421 1550 427
rect 1611 418 1615 428
rect 1371 404 1381 408
rect 1455 406 1460 413
rect 1294 394 1299 403
rect 1377 400 1381 404
rect 1340 397 1381 400
rect 1340 394 1343 397
rect 1377 394 1381 397
rect 1467 406 1472 413
rect 1517 406 1522 416
rect 1567 413 1615 418
rect 1635 427 1841 429
rect 1635 421 1640 427
rect 1672 421 1677 427
rect 1680 426 1841 427
rect 1681 421 1686 426
rect 1832 425 1841 426
rect 1591 406 1596 413
rect 1517 402 1527 406
rect 1276 390 1299 394
rect 1311 390 1343 394
rect 1294 386 1299 390
rect 1351 389 1353 392
rect 1309 377 1314 381
rect 1351 378 1354 389
rect 1368 386 1371 389
rect 1395 378 1398 392
rect 1440 392 1445 401
rect 1523 398 1527 402
rect 1486 395 1527 398
rect 1486 392 1489 395
rect 1523 392 1527 395
rect 1603 406 1608 413
rect 1653 406 1658 416
rect 1653 402 1663 406
rect 1423 388 1445 392
rect 1457 388 1489 392
rect 1440 384 1445 388
rect 1497 387 1499 390
rect 1281 372 1319 377
rect 1281 352 1290 372
rect 1351 373 1398 378
rect 1455 375 1460 379
rect 1497 376 1500 387
rect 1514 384 1517 387
rect 1541 376 1544 390
rect 1576 392 1581 401
rect 1659 398 1663 402
rect 1622 395 1663 398
rect 1622 392 1625 395
rect 1659 392 1663 395
rect 1564 388 1581 392
rect 1593 388 1625 392
rect 1576 384 1581 388
rect 1633 387 1635 390
rect 1430 374 1465 375
rect 1417 370 1465 374
rect 1360 363 1365 364
rect 1417 369 1436 370
rect 1497 371 1544 376
rect 1591 375 1596 379
rect 1633 376 1636 387
rect 1650 384 1653 387
rect 1677 376 1680 390
rect 1566 370 1601 375
rect 1383 363 1388 364
rect 1419 349 1426 369
rect 1506 361 1511 362
rect 1529 361 1534 362
rect 1566 349 1570 370
rect 1633 371 1680 376
rect 1642 361 1647 362
rect 1665 361 1670 362
rect 1290 345 1570 349
rect 1280 344 1570 345
rect 1289 325 1290 330
rect 1441 325 1446 335
rect 1700 340 1785 341
rect 1647 337 1785 340
rect 1647 336 1704 337
rect 1642 325 1647 335
rect 1282 319 1446 325
rect 1223 299 1360 304
rect 1441 303 1446 319
rect 1223 219 1228 299
rect 1355 297 1360 299
rect 1552 320 1647 325
rect 1288 277 1341 283
rect 1383 283 1500 287
rect 1233 239 1276 244
rect 1257 232 1262 239
rect 1269 232 1274 239
rect 1242 219 1247 227
rect 1223 214 1247 219
rect 1259 214 1262 218
rect 1242 210 1247 214
rect 1257 201 1262 205
rect 1288 202 1293 277
rect 1336 271 1341 277
rect 1419 271 1424 283
rect 1431 271 1436 283
rect 1451 282 1500 283
rect 1455 275 1460 282
rect 1467 275 1472 282
rect 1302 260 1307 266
rect 1302 255 1366 260
rect 1385 260 1390 266
rect 1482 261 1487 270
rect 1372 255 1390 260
rect 1302 232 1307 255
rect 1338 249 1341 252
rect 1333 244 1343 249
rect 1336 232 1341 244
rect 1347 235 1353 244
rect 1385 232 1390 255
rect 1437 254 1441 261
rect 1446 257 1470 261
rect 1482 257 1501 261
rect 1420 249 1441 254
rect 1482 253 1487 257
rect 1467 244 1472 248
rect 1451 239 1492 244
rect 1419 202 1424 227
rect 1430 221 1435 224
rect 1451 202 1456 239
rect 1288 201 1451 202
rect 1236 197 1451 201
rect 1236 196 1293 197
rect 1497 193 1501 257
rect 1310 183 1315 187
rect 1332 188 1501 193
rect 1552 189 1557 320
rect 1561 299 1698 304
rect 1561 219 1566 299
rect 1693 297 1698 299
rect 1834 293 1839 425
rect 1988 382 1992 446
rect 2010 442 2015 446
rect 2048 443 2052 446
rect 2099 449 2104 455
rect 2099 444 2115 449
rect 2182 449 2187 455
rect 2121 444 2187 449
rect 2048 438 2069 443
rect 2025 433 2030 437
rect 2004 428 2039 433
rect 2033 391 2038 428
rect 2099 421 2104 444
rect 2148 438 2151 441
rect 2142 433 2156 438
rect 2054 410 2059 413
rect 2133 420 2139 433
rect 2065 391 2070 416
rect 2148 421 2153 433
rect 2182 421 2187 444
rect 2196 391 2201 466
rect 2213 428 2256 433
rect 2215 421 2220 428
rect 2227 421 2232 428
rect 2242 408 2247 416
rect 2261 408 2266 488
rect 2227 403 2230 407
rect 2242 403 2266 408
rect 2242 399 2247 403
rect 2033 390 2201 391
rect 2227 390 2232 394
rect 2033 386 2257 390
rect 2196 385 2257 386
rect 1988 377 2157 382
rect 2152 372 2157 377
rect 2174 372 2179 376
rect 2152 367 2179 372
rect 2117 316 2254 321
rect 2117 314 2122 316
rect 1989 300 2094 304
rect 1989 299 2037 300
rect 1834 287 1907 293
rect 2013 292 2018 299
rect 1626 277 1679 283
rect 1721 283 1907 287
rect 1571 239 1614 244
rect 1595 232 1600 239
rect 1607 232 1612 239
rect 1580 219 1585 227
rect 1561 214 1585 219
rect 1597 214 1600 218
rect 1580 210 1585 214
rect 1595 201 1600 205
rect 1626 202 1631 277
rect 1674 271 1679 277
rect 1757 271 1762 283
rect 1769 271 1774 283
rect 1784 282 1907 283
rect 1787 275 1792 282
rect 1799 275 1804 282
rect 1835 281 1907 282
rect 1640 260 1645 266
rect 1723 260 1728 266
rect 1814 261 1819 270
rect 1640 255 1706 260
rect 1711 255 1728 260
rect 1640 232 1645 255
rect 1676 249 1679 252
rect 1671 244 1689 249
rect 1674 232 1679 244
rect 1689 231 1694 244
rect 1723 232 1728 255
rect 1775 254 1779 261
rect 1784 257 1802 261
rect 1814 257 1839 261
rect 1758 249 1779 254
rect 1814 253 1819 257
rect 1799 244 1804 248
rect 1789 239 1829 244
rect 1757 202 1762 227
rect 1768 221 1773 224
rect 1789 202 1794 239
rect 1626 201 1794 202
rect 1577 197 1794 201
rect 1577 196 1631 197
rect 1835 193 1839 257
rect 1332 183 1337 188
rect 1310 178 1337 183
rect 1552 184 1608 189
rect 1366 152 1372 179
rect 1648 183 1653 187
rect 1670 188 1839 193
rect 1670 183 1675 188
rect 1648 178 1675 183
rect 1547 165 1553 168
rect 1706 165 1711 180
rect 1547 162 1711 165
rect 1893 115 1907 281
rect 2041 288 2046 300
rect 1998 278 2003 287
rect 2053 288 2058 300
rect 2136 294 2189 300
rect 2136 288 2141 294
rect 1976 274 2003 278
rect 2015 274 2027 278
rect 2032 274 2040 278
rect 1976 210 1980 274
rect 1998 270 2003 274
rect 2036 271 2040 274
rect 2087 277 2092 283
rect 2087 272 2102 277
rect 2170 277 2175 283
rect 2109 272 2175 277
rect 2036 266 2057 271
rect 2013 261 2018 265
rect 1993 256 2027 261
rect 2021 219 2026 256
rect 2087 249 2092 272
rect 2136 266 2139 269
rect 2128 261 2144 266
rect 2042 238 2047 241
rect 2121 247 2126 261
rect 2053 219 2058 244
rect 2136 249 2141 261
rect 2170 249 2175 272
rect 2184 219 2189 294
rect 2201 256 2244 261
rect 2203 249 2208 256
rect 2215 249 2220 256
rect 2230 236 2235 244
rect 2249 236 2254 316
rect 2215 231 2218 235
rect 2230 231 2254 236
rect 2230 227 2235 231
rect 2021 218 2189 219
rect 2215 218 2220 222
rect 2021 214 2245 218
rect 2184 213 2245 214
rect 1976 205 2145 210
rect 2140 200 2145 205
rect 2162 200 2167 204
rect 2140 195 2167 200
rect 2108 132 2245 137
rect 2108 130 2113 132
rect 1882 106 1907 115
rect 1978 116 2085 120
rect 1978 115 2028 116
rect 1978 114 1988 115
rect 2004 108 2009 115
rect 1882 105 1901 106
rect 1561 32 1569 36
rect 1427 27 1569 32
rect 1451 20 1456 27
rect 1463 20 1468 27
rect 1490 16 1495 27
rect 1547 16 1552 27
rect 1436 6 1441 15
rect 1184 2 1441 6
rect 1453 2 1479 6
rect 1436 -2 1441 2
rect 1156 -11 1438 -10
rect 1451 -11 1456 -7
rect 1476 -11 1479 2
rect 1499 -11 1504 11
rect 1156 -14 1473 -11
rect 1156 -448 1163 -14
rect 1426 -16 1473 -14
rect 1476 -15 1536 -11
rect 1468 -28 1473 -16
rect 1499 -20 1504 -15
rect 1531 -20 1536 -15
rect 1515 -28 1520 -25
rect 1468 -29 1520 -28
rect 1547 -28 1552 -25
rect 1468 -32 1547 -29
rect 1507 -44 1512 -43
rect 1523 -45 1528 -43
rect 1539 -45 1544 -43
rect 1296 -87 1324 -86
rect 1296 -88 1372 -87
rect 1296 -89 1470 -88
rect 1563 -89 1569 27
rect 1883 -86 1895 105
rect 2032 104 2037 116
rect 1989 94 1994 103
rect 2044 104 2049 116
rect 2127 110 2180 116
rect 2127 104 2132 110
rect 1967 90 1994 94
rect 2006 90 2018 94
rect 2023 90 2031 94
rect 1967 26 1971 90
rect 1989 86 1994 90
rect 2027 87 2031 90
rect 2078 93 2083 99
rect 2078 88 2094 93
rect 2161 93 2166 99
rect 2100 88 2166 93
rect 2027 82 2048 87
rect 2004 77 2009 81
rect 1984 72 2018 77
rect 2012 35 2017 72
rect 2078 65 2083 88
rect 2127 82 2130 85
rect 2119 77 2135 82
rect 2033 54 2038 57
rect 2112 67 2117 77
rect 2127 65 2132 77
rect 2161 65 2166 88
rect 2044 35 2049 60
rect 2175 35 2180 110
rect 2192 72 2235 77
rect 2194 65 2199 72
rect 2206 65 2211 72
rect 2221 52 2226 60
rect 2240 52 2245 132
rect 2206 47 2209 51
rect 2221 47 2245 52
rect 2221 43 2226 47
rect 2012 34 2180 35
rect 2206 34 2211 38
rect 2012 30 2236 34
rect 2175 29 2236 30
rect 1967 25 1976 26
rect 1984 25 2136 26
rect 1967 22 2136 25
rect 1967 21 1976 22
rect 1984 21 2136 22
rect 2131 16 2136 21
rect 2153 16 2158 20
rect 2131 11 2158 16
rect 1575 -89 1606 -88
rect 1800 -89 1895 -86
rect 1296 -90 1895 -89
rect 1297 -101 1301 -90
rect 1227 -105 1301 -101
rect 1321 -92 1895 -90
rect 1321 -98 1326 -92
rect 1358 -98 1363 -92
rect 1367 -98 1372 -92
rect 1443 -103 1447 -92
rect 1173 -139 1207 -136
rect 1173 -445 1176 -139
rect 1202 -190 1207 -139
rect 1227 -205 1233 -105
rect 1253 -106 1301 -105
rect 1277 -113 1282 -106
rect 1289 -113 1294 -106
rect 1339 -113 1344 -103
rect 1399 -108 1447 -103
rect 1467 -93 1583 -92
rect 1467 -94 1518 -93
rect 1467 -100 1472 -94
rect 1504 -100 1509 -94
rect 1513 -100 1518 -94
rect 1579 -103 1583 -93
rect 1339 -117 1349 -113
rect 1423 -115 1428 -108
rect 1262 -127 1267 -118
rect 1345 -121 1349 -117
rect 1308 -124 1349 -121
rect 1308 -127 1311 -124
rect 1345 -127 1349 -124
rect 1435 -115 1440 -108
rect 1485 -115 1490 -105
rect 1535 -108 1583 -103
rect 1603 -94 1895 -92
rect 1603 -100 1608 -94
rect 1640 -100 1645 -94
rect 1648 -95 1895 -94
rect 1649 -100 1654 -95
rect 1559 -115 1564 -108
rect 1485 -119 1495 -115
rect 1244 -131 1267 -127
rect 1279 -131 1311 -127
rect 1262 -135 1267 -131
rect 1319 -132 1321 -129
rect 1277 -144 1282 -140
rect 1319 -143 1322 -132
rect 1336 -135 1339 -132
rect 1363 -143 1366 -129
rect 1408 -129 1413 -120
rect 1491 -123 1495 -119
rect 1454 -126 1495 -123
rect 1454 -129 1457 -126
rect 1491 -129 1495 -126
rect 1571 -115 1576 -108
rect 1621 -115 1626 -105
rect 1621 -119 1631 -115
rect 1391 -133 1413 -129
rect 1425 -133 1457 -129
rect 1408 -137 1413 -133
rect 1465 -134 1467 -131
rect 1249 -149 1287 -144
rect 1249 -169 1258 -149
rect 1319 -148 1366 -143
rect 1423 -146 1428 -142
rect 1465 -145 1468 -134
rect 1482 -137 1485 -134
rect 1509 -145 1512 -131
rect 1544 -129 1549 -120
rect 1627 -123 1631 -119
rect 1590 -126 1631 -123
rect 1590 -129 1593 -126
rect 1627 -129 1631 -126
rect 1532 -133 1549 -129
rect 1561 -133 1593 -129
rect 1544 -137 1549 -133
rect 1601 -134 1603 -131
rect 1398 -147 1433 -146
rect 1385 -151 1433 -147
rect 1328 -158 1333 -157
rect 1385 -152 1404 -151
rect 1465 -150 1512 -145
rect 1559 -146 1564 -142
rect 1601 -145 1604 -134
rect 1618 -137 1621 -134
rect 1645 -145 1648 -131
rect 1534 -151 1569 -146
rect 1351 -158 1356 -157
rect 1387 -172 1394 -152
rect 1474 -160 1479 -159
rect 1497 -160 1502 -159
rect 1534 -172 1538 -151
rect 1601 -150 1648 -145
rect 1610 -160 1615 -159
rect 1633 -160 1638 -159
rect 1258 -176 1538 -172
rect 1248 -177 1538 -176
rect 1257 -196 1258 -191
rect 1409 -196 1414 -186
rect 1668 -181 1753 -180
rect 1615 -184 1753 -181
rect 1615 -185 1672 -184
rect 1610 -196 1615 -186
rect 1250 -202 1414 -196
rect 1191 -222 1328 -217
rect 1409 -218 1414 -202
rect 1191 -302 1196 -222
rect 1323 -224 1328 -222
rect 1520 -201 1615 -196
rect 1256 -244 1309 -238
rect 1351 -238 1468 -234
rect 1201 -282 1244 -277
rect 1225 -289 1230 -282
rect 1237 -289 1242 -282
rect 1210 -302 1215 -294
rect 1191 -307 1215 -302
rect 1227 -307 1230 -303
rect 1210 -311 1215 -307
rect 1225 -320 1230 -316
rect 1256 -319 1261 -244
rect 1304 -250 1309 -244
rect 1387 -250 1392 -238
rect 1399 -250 1404 -238
rect 1419 -239 1468 -238
rect 1423 -246 1428 -239
rect 1435 -246 1440 -239
rect 1270 -261 1275 -255
rect 1270 -266 1334 -261
rect 1353 -261 1358 -255
rect 1450 -260 1455 -251
rect 1340 -266 1358 -261
rect 1270 -289 1275 -266
rect 1306 -272 1309 -269
rect 1301 -277 1319 -272
rect 1304 -289 1309 -277
rect 1319 -291 1324 -277
rect 1353 -289 1358 -266
rect 1405 -267 1409 -260
rect 1414 -264 1438 -260
rect 1450 -264 1469 -260
rect 1388 -272 1409 -267
rect 1450 -268 1455 -264
rect 1435 -277 1440 -273
rect 1419 -282 1460 -277
rect 1387 -319 1392 -294
rect 1398 -300 1403 -297
rect 1419 -319 1424 -282
rect 1256 -320 1419 -319
rect 1204 -324 1419 -320
rect 1204 -325 1261 -324
rect 1465 -328 1469 -264
rect 1278 -338 1283 -334
rect 1300 -333 1469 -328
rect 1520 -332 1525 -201
rect 1529 -222 1666 -217
rect 1529 -302 1534 -222
rect 1661 -224 1666 -222
rect 1802 -234 1807 -95
rect 1883 -97 1895 -95
rect 1828 -234 1833 -232
rect 1594 -244 1647 -238
rect 1689 -238 1833 -234
rect 1539 -282 1582 -277
rect 1563 -289 1568 -282
rect 1575 -289 1580 -282
rect 1548 -302 1553 -294
rect 1529 -307 1553 -302
rect 1565 -307 1568 -303
rect 1548 -311 1553 -307
rect 1563 -320 1568 -316
rect 1594 -319 1599 -244
rect 1642 -250 1647 -244
rect 1725 -250 1730 -238
rect 1737 -250 1742 -238
rect 1752 -239 1833 -238
rect 1755 -246 1760 -239
rect 1767 -246 1772 -239
rect 1608 -261 1613 -255
rect 1691 -261 1696 -255
rect 1782 -260 1787 -251
rect 1608 -266 1674 -261
rect 1679 -266 1696 -261
rect 1608 -289 1613 -266
rect 1644 -272 1647 -269
rect 1639 -277 1657 -272
rect 1642 -289 1647 -277
rect 1657 -290 1663 -278
rect 1691 -289 1696 -266
rect 1743 -267 1747 -260
rect 1752 -264 1770 -260
rect 1782 -264 1807 -260
rect 1726 -272 1747 -267
rect 1782 -268 1787 -264
rect 1767 -277 1772 -273
rect 1757 -282 1797 -277
rect 1725 -319 1730 -294
rect 1736 -300 1741 -297
rect 1757 -319 1762 -282
rect 1594 -320 1762 -319
rect 1545 -324 1762 -320
rect 1545 -325 1599 -324
rect 1803 -328 1807 -264
rect 1300 -338 1305 -333
rect 1278 -343 1305 -338
rect 1520 -337 1576 -332
rect 1334 -358 1340 -342
rect 1616 -338 1621 -334
rect 1638 -333 1807 -328
rect 1638 -338 1643 -333
rect 1616 -343 1643 -338
rect 1515 -356 1521 -353
rect 1674 -356 1679 -341
rect 1515 -359 1679 -356
rect 1427 -424 1569 -419
rect 1451 -431 1456 -424
rect 1463 -431 1468 -424
rect 1490 -435 1495 -424
rect 1547 -435 1552 -424
rect 1436 -445 1441 -436
rect 1173 -448 1441 -445
rect 1157 -463 1163 -448
rect 1351 -449 1441 -448
rect 1453 -449 1479 -445
rect 1436 -453 1441 -449
rect 1451 -462 1456 -458
rect 1476 -462 1479 -449
rect 1499 -462 1504 -440
rect 1426 -463 1473 -462
rect 1157 -467 1473 -463
rect 1476 -466 1536 -462
rect 1157 -481 1163 -467
rect 1156 -912 1163 -481
rect 1468 -479 1473 -467
rect 1499 -471 1504 -466
rect 1531 -471 1536 -466
rect 1515 -479 1520 -476
rect 1468 -480 1520 -479
rect 1547 -479 1552 -476
rect 1468 -483 1547 -480
rect 1507 -495 1512 -494
rect 1523 -496 1528 -494
rect 1539 -496 1544 -494
rect 1296 -538 1324 -537
rect 1296 -539 1372 -538
rect 1296 -540 1470 -539
rect 1563 -540 1569 -424
rect 1575 -540 1606 -539
rect 1802 -540 1807 -539
rect 1296 -541 1807 -540
rect 1828 -541 1833 -239
rect 1297 -552 1301 -541
rect 1227 -556 1301 -552
rect 1321 -543 1833 -541
rect 1321 -549 1326 -543
rect 1358 -549 1363 -543
rect 1367 -549 1372 -543
rect 1443 -554 1447 -543
rect 1171 -592 1207 -586
rect 1171 -871 1174 -592
rect 1202 -641 1207 -592
rect 1227 -656 1233 -556
rect 1253 -557 1301 -556
rect 1277 -564 1282 -557
rect 1289 -564 1294 -557
rect 1339 -564 1344 -554
rect 1399 -559 1447 -554
rect 1467 -544 1583 -543
rect 1467 -545 1518 -544
rect 1467 -551 1472 -545
rect 1504 -551 1509 -545
rect 1513 -551 1518 -545
rect 1579 -554 1583 -544
rect 1339 -568 1349 -564
rect 1423 -566 1428 -559
rect 1262 -578 1267 -569
rect 1345 -572 1349 -568
rect 1308 -575 1349 -572
rect 1308 -578 1311 -575
rect 1345 -578 1349 -575
rect 1435 -566 1440 -559
rect 1485 -566 1490 -556
rect 1535 -559 1583 -554
rect 1603 -545 1833 -543
rect 1603 -551 1608 -545
rect 1640 -551 1645 -545
rect 1648 -546 1807 -545
rect 1649 -551 1654 -546
rect 1559 -566 1564 -559
rect 1485 -570 1495 -566
rect 1244 -582 1267 -578
rect 1279 -582 1311 -578
rect 1262 -586 1267 -582
rect 1319 -583 1321 -580
rect 1277 -595 1282 -591
rect 1319 -594 1322 -583
rect 1336 -586 1339 -583
rect 1363 -594 1366 -580
rect 1408 -580 1413 -571
rect 1491 -574 1495 -570
rect 1454 -577 1495 -574
rect 1454 -580 1457 -577
rect 1491 -580 1495 -577
rect 1571 -566 1576 -559
rect 1621 -566 1626 -556
rect 1621 -570 1631 -566
rect 1391 -584 1413 -580
rect 1425 -584 1457 -580
rect 1408 -588 1413 -584
rect 1465 -585 1467 -582
rect 1249 -600 1287 -595
rect 1249 -620 1258 -600
rect 1319 -599 1366 -594
rect 1423 -597 1428 -593
rect 1465 -596 1468 -585
rect 1482 -588 1485 -585
rect 1509 -596 1512 -582
rect 1544 -580 1549 -571
rect 1627 -574 1631 -570
rect 1590 -577 1631 -574
rect 1590 -580 1593 -577
rect 1627 -580 1631 -577
rect 1532 -584 1549 -580
rect 1561 -584 1593 -580
rect 1544 -588 1549 -584
rect 1601 -585 1603 -582
rect 1398 -598 1433 -597
rect 1385 -602 1433 -598
rect 1328 -609 1333 -608
rect 1385 -603 1404 -602
rect 1465 -601 1512 -596
rect 1559 -597 1564 -593
rect 1601 -596 1604 -585
rect 1618 -588 1621 -585
rect 1645 -596 1648 -582
rect 1534 -602 1569 -597
rect 1351 -609 1356 -608
rect 1387 -623 1394 -603
rect 1474 -611 1479 -610
rect 1497 -611 1502 -610
rect 1534 -623 1538 -602
rect 1601 -601 1648 -596
rect 1610 -611 1615 -610
rect 1633 -611 1638 -610
rect 1258 -627 1538 -623
rect 1248 -628 1538 -627
rect 1257 -647 1258 -642
rect 1409 -647 1414 -637
rect 1668 -632 1753 -631
rect 1615 -635 1753 -632
rect 1615 -636 1672 -635
rect 1610 -647 1615 -637
rect 1250 -653 1414 -647
rect 1191 -673 1328 -668
rect 1409 -669 1414 -653
rect 1191 -753 1196 -673
rect 1323 -675 1328 -673
rect 1520 -652 1615 -647
rect 1256 -695 1309 -689
rect 1351 -689 1468 -685
rect 1201 -733 1244 -728
rect 1225 -740 1230 -733
rect 1237 -740 1242 -733
rect 1210 -753 1215 -745
rect 1191 -758 1215 -753
rect 1227 -758 1230 -754
rect 1210 -762 1215 -758
rect 1225 -771 1230 -767
rect 1256 -770 1261 -695
rect 1304 -701 1309 -695
rect 1387 -701 1392 -689
rect 1399 -701 1404 -689
rect 1419 -690 1468 -689
rect 1423 -697 1428 -690
rect 1435 -697 1440 -690
rect 1270 -712 1275 -706
rect 1270 -717 1334 -712
rect 1353 -712 1358 -706
rect 1450 -711 1455 -702
rect 1340 -717 1358 -712
rect 1270 -740 1275 -717
rect 1306 -723 1309 -720
rect 1301 -728 1319 -723
rect 1304 -740 1309 -728
rect 1319 -742 1324 -728
rect 1353 -740 1358 -717
rect 1405 -718 1409 -711
rect 1414 -715 1438 -711
rect 1450 -715 1469 -711
rect 1388 -723 1409 -718
rect 1450 -719 1455 -715
rect 1435 -728 1440 -724
rect 1419 -733 1460 -728
rect 1387 -770 1392 -745
rect 1398 -751 1403 -748
rect 1419 -770 1424 -733
rect 1256 -771 1419 -770
rect 1204 -775 1419 -771
rect 1204 -776 1261 -775
rect 1465 -779 1469 -715
rect 1278 -789 1283 -785
rect 1300 -784 1469 -779
rect 1520 -783 1525 -652
rect 1529 -673 1666 -668
rect 1529 -753 1534 -673
rect 1661 -675 1666 -673
rect 1802 -674 1807 -546
rect 1802 -678 1827 -674
rect 1802 -685 1807 -678
rect 1594 -695 1647 -689
rect 1689 -689 1807 -685
rect 1539 -733 1582 -728
rect 1563 -740 1568 -733
rect 1575 -740 1580 -733
rect 1548 -753 1553 -745
rect 1529 -758 1553 -753
rect 1565 -758 1568 -754
rect 1548 -762 1553 -758
rect 1563 -771 1568 -767
rect 1594 -770 1599 -695
rect 1642 -701 1647 -695
rect 1725 -701 1730 -689
rect 1737 -701 1742 -689
rect 1752 -690 1807 -689
rect 1755 -697 1760 -690
rect 1767 -697 1772 -690
rect 1608 -712 1613 -706
rect 1691 -712 1696 -706
rect 1782 -711 1787 -702
rect 1608 -717 1674 -712
rect 1679 -717 1696 -712
rect 1608 -740 1613 -717
rect 1644 -723 1647 -720
rect 1639 -728 1659 -723
rect 1642 -740 1647 -728
rect 1655 -738 1661 -728
rect 1691 -740 1696 -717
rect 1743 -718 1747 -711
rect 1752 -715 1770 -711
rect 1782 -715 1807 -711
rect 1726 -723 1747 -718
rect 1782 -719 1787 -715
rect 1767 -728 1772 -724
rect 1757 -733 1797 -728
rect 1725 -770 1730 -745
rect 1736 -751 1741 -748
rect 1757 -770 1762 -733
rect 1594 -771 1762 -770
rect 1545 -775 1762 -771
rect 1545 -776 1599 -775
rect 1803 -779 1807 -715
rect 1300 -789 1305 -784
rect 1278 -794 1305 -789
rect 1520 -788 1576 -783
rect 1334 -809 1340 -793
rect 1616 -789 1621 -785
rect 1638 -784 1807 -779
rect 1638 -789 1643 -784
rect 1616 -794 1643 -789
rect 1515 -807 1521 -804
rect 1674 -807 1679 -792
rect 1515 -810 1679 -807
rect 1171 -874 1385 -871
rect 1418 -874 1554 -869
rect 1381 -895 1385 -874
rect 1442 -881 1447 -874
rect 1454 -881 1459 -874
rect 1481 -885 1486 -874
rect 1538 -885 1543 -874
rect 1427 -895 1432 -886
rect 1381 -899 1432 -895
rect 1444 -899 1470 -895
rect 1427 -903 1432 -899
rect 1442 -912 1447 -908
rect 1467 -912 1470 -899
rect 1490 -912 1495 -890
rect 1154 -916 1464 -912
rect 1467 -916 1527 -912
rect 1417 -917 1464 -916
rect 1459 -929 1464 -917
rect 1490 -921 1495 -916
rect 1522 -921 1527 -916
rect 1506 -929 1511 -926
rect 1459 -930 1511 -929
rect 1538 -929 1543 -926
rect 1459 -933 1538 -930
rect 1498 -945 1503 -944
rect 1514 -946 1519 -944
rect 1530 -946 1535 -944
rect 1287 -988 1315 -987
rect 1287 -989 1363 -988
rect 1287 -990 1461 -989
rect 1554 -990 1560 -876
rect 1566 -990 1597 -989
rect 1793 -990 1798 -989
rect 1822 -990 1827 -678
rect 1287 -991 1798 -990
rect 1806 -991 1827 -990
rect 1288 -1002 1292 -991
rect 1218 -1006 1292 -1002
rect 1312 -993 1827 -991
rect 1312 -999 1317 -993
rect 1349 -999 1354 -993
rect 1358 -999 1363 -993
rect 1434 -1004 1438 -993
rect 1193 -1091 1198 -1042
rect 1218 -1106 1224 -1006
rect 1244 -1007 1292 -1006
rect 1268 -1014 1273 -1007
rect 1280 -1014 1285 -1007
rect 1330 -1014 1335 -1004
rect 1390 -1009 1438 -1004
rect 1458 -994 1574 -993
rect 1458 -995 1509 -994
rect 1458 -1001 1463 -995
rect 1495 -1001 1500 -995
rect 1504 -1001 1509 -995
rect 1570 -1004 1574 -994
rect 1330 -1018 1340 -1014
rect 1414 -1016 1419 -1009
rect 1253 -1028 1258 -1019
rect 1336 -1022 1340 -1018
rect 1299 -1025 1340 -1022
rect 1299 -1028 1302 -1025
rect 1336 -1028 1340 -1025
rect 1426 -1016 1431 -1009
rect 1476 -1016 1481 -1006
rect 1526 -1009 1574 -1004
rect 1594 -995 1827 -993
rect 1594 -1001 1599 -995
rect 1631 -1001 1636 -995
rect 1639 -996 1817 -995
rect 1640 -1001 1645 -996
rect 1550 -1016 1555 -1009
rect 1476 -1020 1486 -1016
rect 1235 -1032 1258 -1028
rect 1270 -1032 1302 -1028
rect 1253 -1036 1258 -1032
rect 1310 -1033 1312 -1030
rect 1268 -1045 1273 -1041
rect 1310 -1044 1313 -1033
rect 1327 -1036 1330 -1033
rect 1354 -1044 1357 -1030
rect 1399 -1030 1404 -1021
rect 1482 -1024 1486 -1020
rect 1445 -1027 1486 -1024
rect 1445 -1030 1448 -1027
rect 1482 -1030 1486 -1027
rect 1562 -1016 1567 -1009
rect 1612 -1016 1617 -1006
rect 1612 -1020 1622 -1016
rect 1382 -1034 1404 -1030
rect 1416 -1034 1448 -1030
rect 1399 -1038 1404 -1034
rect 1456 -1035 1458 -1032
rect 1240 -1050 1278 -1045
rect 1240 -1070 1249 -1050
rect 1310 -1049 1357 -1044
rect 1414 -1047 1419 -1043
rect 1456 -1046 1459 -1035
rect 1473 -1038 1476 -1035
rect 1500 -1046 1503 -1032
rect 1535 -1030 1540 -1021
rect 1618 -1024 1622 -1020
rect 1581 -1027 1622 -1024
rect 1581 -1030 1584 -1027
rect 1618 -1030 1622 -1027
rect 1523 -1034 1540 -1030
rect 1552 -1034 1584 -1030
rect 1535 -1038 1540 -1034
rect 1592 -1035 1594 -1032
rect 1389 -1048 1424 -1047
rect 1376 -1052 1424 -1048
rect 1319 -1059 1324 -1058
rect 1376 -1053 1395 -1052
rect 1456 -1051 1503 -1046
rect 1550 -1047 1555 -1043
rect 1592 -1046 1595 -1035
rect 1609 -1038 1612 -1035
rect 1636 -1046 1639 -1032
rect 1525 -1052 1560 -1047
rect 1342 -1059 1347 -1058
rect 1378 -1073 1385 -1053
rect 1465 -1061 1470 -1060
rect 1488 -1061 1493 -1060
rect 1525 -1073 1529 -1052
rect 1592 -1051 1639 -1046
rect 1601 -1061 1606 -1060
rect 1624 -1061 1629 -1060
rect 1249 -1077 1529 -1073
rect 1239 -1078 1529 -1077
rect 1248 -1097 1249 -1092
rect 1400 -1097 1405 -1087
rect 1659 -1082 1744 -1081
rect 1606 -1085 1744 -1082
rect 1606 -1086 1663 -1085
rect 1601 -1097 1606 -1087
rect 1241 -1103 1405 -1097
rect 1219 -1115 1224 -1114
rect 1182 -1123 1319 -1118
rect 1400 -1119 1405 -1103
rect 1182 -1203 1187 -1123
rect 1314 -1125 1319 -1123
rect 1511 -1102 1606 -1097
rect 1247 -1145 1300 -1139
rect 1342 -1139 1459 -1135
rect 1192 -1183 1235 -1178
rect 1216 -1190 1221 -1183
rect 1228 -1190 1233 -1183
rect 1201 -1203 1206 -1195
rect 1182 -1208 1206 -1203
rect 1218 -1208 1221 -1204
rect 1201 -1212 1206 -1208
rect 1216 -1221 1221 -1217
rect 1247 -1220 1252 -1145
rect 1295 -1151 1300 -1145
rect 1378 -1151 1383 -1139
rect 1390 -1151 1395 -1139
rect 1410 -1140 1459 -1139
rect 1414 -1147 1419 -1140
rect 1426 -1147 1431 -1140
rect 1261 -1162 1266 -1156
rect 1344 -1162 1349 -1156
rect 1441 -1161 1446 -1152
rect 1261 -1167 1349 -1162
rect 1261 -1190 1266 -1167
rect 1292 -1178 1312 -1173
rect 1295 -1190 1300 -1178
rect 1308 -1190 1312 -1178
rect 1344 -1190 1349 -1167
rect 1396 -1168 1400 -1161
rect 1405 -1165 1429 -1161
rect 1441 -1165 1460 -1161
rect 1379 -1173 1400 -1168
rect 1441 -1169 1446 -1165
rect 1426 -1178 1431 -1174
rect 1410 -1183 1451 -1178
rect 1378 -1220 1383 -1195
rect 1389 -1201 1394 -1198
rect 1410 -1220 1415 -1183
rect 1247 -1221 1410 -1220
rect 1195 -1225 1410 -1221
rect 1195 -1226 1252 -1225
rect 1456 -1229 1460 -1165
rect 1269 -1239 1274 -1235
rect 1291 -1234 1460 -1229
rect 1511 -1233 1516 -1102
rect 1520 -1123 1657 -1118
rect 1520 -1203 1525 -1123
rect 1652 -1125 1657 -1123
rect 1793 -1135 1798 -996
rect 1585 -1145 1638 -1139
rect 1680 -1139 1798 -1135
rect 1530 -1183 1573 -1178
rect 1554 -1190 1559 -1183
rect 1566 -1190 1571 -1183
rect 1539 -1203 1544 -1195
rect 1520 -1208 1544 -1203
rect 1556 -1208 1559 -1204
rect 1539 -1212 1544 -1208
rect 1554 -1221 1559 -1217
rect 1585 -1220 1590 -1145
rect 1633 -1151 1638 -1145
rect 1716 -1151 1721 -1139
rect 1728 -1151 1733 -1139
rect 1743 -1140 1798 -1139
rect 1746 -1147 1751 -1140
rect 1758 -1147 1763 -1140
rect 1599 -1162 1604 -1156
rect 1682 -1162 1687 -1156
rect 1773 -1161 1778 -1152
rect 1599 -1167 1665 -1162
rect 1670 -1167 1687 -1162
rect 1599 -1190 1604 -1167
rect 1630 -1178 1648 -1173
rect 1633 -1190 1638 -1178
rect 1648 -1192 1653 -1178
rect 1682 -1190 1687 -1167
rect 1734 -1168 1738 -1161
rect 1743 -1165 1761 -1161
rect 1773 -1165 1798 -1161
rect 1717 -1173 1738 -1168
rect 1773 -1169 1778 -1165
rect 1758 -1178 1763 -1174
rect 1748 -1183 1788 -1178
rect 1716 -1220 1721 -1195
rect 1727 -1201 1732 -1198
rect 1748 -1220 1753 -1183
rect 1585 -1221 1753 -1220
rect 1536 -1225 1753 -1221
rect 1536 -1226 1590 -1225
rect 1794 -1229 1798 -1165
rect 1291 -1239 1296 -1234
rect 1511 -1238 1567 -1233
rect 1269 -1244 1296 -1239
rect 1607 -1239 1612 -1235
rect 1629 -1234 1798 -1229
rect 1629 -1239 1634 -1234
rect 1607 -1244 1634 -1239
rect 1506 -1257 1512 -1254
rect 1665 -1257 1670 -1242
rect 1506 -1260 1670 -1257
<< m2contact >>
rect 944 1553 949 1558
rect 895 1543 902 1550
rect 936 1528 941 1535
rect 859 1517 869 1522
rect 944 1517 950 1522
rect 943 1493 949 1499
rect 882 1462 889 1469
rect 669 1426 674 1433
rect 866 1430 872 1439
rect 700 1424 707 1430
rect 795 1413 800 1419
rect 132 1335 141 1346
rect 655 1397 661 1402
rect 795 1397 802 1402
rect 1071 1386 1086 1395
rect 655 1377 662 1382
rect 795 1377 802 1382
rect 931 1379 936 1384
rect 186 1310 199 1320
rect 75 1296 86 1306
rect 461 1294 475 1304
rect 186 1266 193 1272
rect 229 1241 234 1246
rect 356 1266 361 1271
rect 227 1223 232 1228
rect 287 1240 294 1245
rect 250 1223 255 1228
rect 304 1200 309 1205
rect 383 1228 390 1235
rect 398 1226 403 1233
rect 458 1223 463 1228
rect 530 1282 538 1290
rect 604 1356 615 1363
rect 655 1356 663 1362
rect 736 1357 750 1362
rect 795 1359 802 1364
rect 578 1234 587 1248
rect 931 1358 937 1363
rect 840 1322 853 1338
rect 655 1312 664 1319
rect 681 1310 690 1318
rect 796 1315 801 1321
rect 899 1322 909 1331
rect 1077 1325 1088 1336
rect 1176 1319 1187 1328
rect 2362 1355 2371 1364
rect 2071 1340 2083 1351
rect 796 1291 801 1298
rect 615 1276 622 1281
rect 961 1275 967 1283
rect 1116 1258 1126 1264
rect 1206 1250 1211 1255
rect 1157 1240 1164 1247
rect 690 1229 695 1235
rect 706 1229 711 1235
rect 754 1229 759 1236
rect 472 1198 477 1203
rect 720 1199 730 1207
rect 755 1205 765 1213
rect 545 1181 561 1193
rect 503 1132 517 1141
rect 224 1072 229 1077
rect 183 1043 190 1049
rect 226 1019 231 1024
rect 353 1044 358 1049
rect 224 1001 229 1006
rect 286 1015 292 1021
rect 247 1001 252 1006
rect 379 1006 388 1011
rect 301 978 306 983
rect 455 1001 460 1006
rect 469 976 474 981
rect 568 1180 585 1191
rect 548 1131 560 1143
rect 621 1156 633 1167
rect 570 1114 581 1129
rect 541 1091 552 1102
rect 739 1175 751 1191
rect 914 1162 925 1171
rect 1198 1225 1203 1232
rect 1221 1225 1226 1232
rect 1012 1156 1024 1163
rect 1039 1156 1051 1163
rect 779 1112 789 1119
rect 815 1110 828 1120
rect 716 1095 727 1106
rect 958 1093 970 1107
rect 1102 1101 1117 1110
rect 1318 1087 1326 1094
rect 573 1064 585 1074
rect 651 1065 662 1074
rect 1663 1295 1676 1308
rect 1991 1296 1998 1304
rect 2618 1327 2628 1336
rect 2186 1311 2194 1318
rect 2114 1303 2124 1310
rect 2132 1291 2142 1299
rect 2262 1307 2271 1313
rect 2766 1304 2776 1314
rect 2281 1292 2289 1298
rect 1887 1224 1892 1229
rect 1980 1231 1986 1238
rect 1934 1214 1941 1221
rect 2023 1224 2028 1229
rect 2118 1232 2124 1239
rect 1872 1199 1877 1206
rect 1895 1199 1900 1206
rect 2070 1214 2077 1221
rect 2169 1226 2174 1231
rect 2264 1233 2270 1240
rect 2216 1216 2223 1223
rect 2316 1226 2321 1231
rect 2420 1233 2427 1241
rect 2008 1199 2013 1206
rect 2031 1199 2036 1206
rect 2154 1201 2159 1208
rect 2177 1201 2182 1208
rect 2363 1216 2370 1223
rect 2528 1225 2533 1230
rect 2281 1200 2289 1206
rect 2301 1201 2306 1208
rect 2324 1201 2329 1208
rect 2575 1215 2582 1222
rect 2664 1225 2669 1230
rect 2513 1200 2518 1207
rect 2536 1200 2541 1207
rect 2711 1215 2718 1222
rect 2810 1227 2815 1232
rect 2857 1217 2864 1224
rect 2957 1227 2962 1232
rect 2649 1200 2654 1207
rect 2672 1200 2677 1207
rect 2795 1202 2800 1209
rect 2818 1202 2823 1209
rect 3004 1217 3011 1224
rect 2942 1202 2947 1209
rect 2965 1202 2970 1209
rect 1887 1116 1892 1121
rect 1993 1124 1998 1130
rect 1934 1106 1941 1113
rect 2031 1116 2036 1121
rect 2133 1122 2139 1129
rect 1832 1086 1838 1093
rect 1872 1090 1877 1098
rect 1895 1091 1900 1098
rect 660 1013 667 1019
rect 759 1004 764 1009
rect 815 1014 821 1019
rect 710 994 717 1001
rect 906 1004 911 1009
rect 959 1011 966 1017
rect 153 933 160 940
rect 198 934 205 941
rect 480 893 489 903
rect 144 881 152 887
rect 45 833 50 838
rect 161 859 168 865
rect 356 859 361 864
rect 228 832 233 838
rect 227 816 232 821
rect 147 800 153 806
rect 186 800 192 805
rect 226 788 231 794
rect 143 776 151 782
rect 288 831 293 836
rect 250 816 255 821
rect 304 793 309 798
rect 383 821 391 826
rect 458 816 463 821
rect 472 791 477 796
rect 542 965 554 976
rect 572 971 583 981
rect 751 979 756 986
rect 774 979 779 986
rect 857 994 864 1001
rect 1052 1002 1057 1007
rect 1103 1009 1109 1014
rect 898 979 903 986
rect 1003 992 1010 999
rect 1188 1002 1193 1007
rect 921 979 926 986
rect 1044 977 1049 984
rect 1067 977 1072 984
rect 1139 992 1146 999
rect 1180 977 1185 984
rect 1203 977 1208 984
rect 541 909 551 922
rect 535 882 545 890
rect 635 906 641 911
rect 620 857 630 867
rect 501 758 510 765
rect 502 729 509 736
rect 510 701 516 709
rect 186 684 193 690
rect 356 684 361 689
rect 228 658 233 663
rect 227 641 232 646
rect 288 656 294 661
rect 250 641 255 646
rect 378 646 388 651
rect 304 618 309 623
rect 458 641 463 646
rect 472 616 477 621
rect 617 628 626 640
rect 476 571 485 581
rect 1580 1046 1585 1051
rect 1660 1055 1666 1060
rect 2078 1106 2085 1113
rect 2180 1118 2185 1123
rect 2282 1125 2288 1131
rect 2227 1108 2234 1115
rect 2325 1119 2330 1124
rect 2407 1125 2415 1132
rect 2372 1109 2379 1116
rect 2016 1091 2021 1098
rect 2039 1091 2044 1098
rect 2165 1093 2170 1100
rect 2188 1093 2193 1100
rect 2310 1093 2315 1100
rect 2333 1094 2338 1101
rect 1627 1037 1634 1043
rect 1488 1015 1496 1023
rect 1565 1022 1570 1029
rect 1656 1034 1665 1043
rect 1832 1051 1838 1056
rect 1588 1023 1593 1029
rect 662 904 668 910
rect 750 897 755 902
rect 804 906 809 911
rect 701 887 708 894
rect 895 896 900 901
rect 945 902 952 907
rect 742 872 747 879
rect 765 871 770 878
rect 846 886 853 893
rect 1044 894 1049 899
rect 1090 903 1095 908
rect 1405 916 1410 921
rect 1429 916 1435 921
rect 1442 916 1447 921
rect 1465 916 1473 921
rect 887 871 892 878
rect 910 871 915 878
rect 995 884 1002 891
rect 1188 894 1193 899
rect 1337 896 1353 908
rect 1036 869 1041 876
rect 1059 869 1064 876
rect 1139 884 1146 891
rect 1180 869 1185 876
rect 1203 868 1208 876
rect 1244 868 1249 874
rect 1318 868 1323 874
rect 1441 894 1447 899
rect 1319 704 1326 710
rect 1720 1036 1729 1045
rect 1791 1018 1796 1023
rect 1666 937 1671 942
rect 1579 928 1584 933
rect 1624 919 1632 924
rect 1564 903 1569 908
rect 1586 902 1592 908
rect 1848 1008 1855 1017
rect 2383 993 2388 998
rect 1732 937 1738 942
rect 2218 927 2223 932
rect 2373 947 2379 952
rect 2288 936 2293 941
rect 2335 926 2342 933
rect 2424 936 2429 941
rect 2506 944 2511 950
rect 2273 911 2278 918
rect 2296 911 2301 918
rect 1762 894 1769 902
rect 2099 884 2104 889
rect 2471 926 2478 933
rect 2648 947 2653 952
rect 2570 938 2575 943
rect 2617 928 2624 935
rect 2717 938 2722 943
rect 2818 946 2825 954
rect 2409 911 2414 918
rect 2432 911 2437 918
rect 2555 913 2560 920
rect 2578 913 2583 920
rect 2764 928 2771 935
rect 2702 913 2707 920
rect 2725 913 2730 920
rect 1670 833 1678 839
rect 1578 824 1583 829
rect 1623 815 1631 821
rect 1545 776 1555 782
rect 2002 761 2007 766
rect 1578 728 1583 733
rect 1805 736 1815 743
rect 1624 718 1632 724
rect 1769 718 1774 723
rect 1586 704 1591 711
rect 1938 717 1944 722
rect 2006 689 2011 694
rect 2288 828 2293 833
rect 2367 837 2372 842
rect 2335 818 2342 825
rect 2520 837 2525 842
rect 2432 828 2437 833
rect 2273 802 2278 810
rect 2296 803 2301 810
rect 2479 818 2486 825
rect 2667 839 2674 844
rect 2581 830 2586 835
rect 2628 820 2635 827
rect 2812 840 2819 845
rect 2726 831 2731 836
rect 2773 821 2780 828
rect 2417 803 2422 810
rect 2440 803 2445 810
rect 2566 805 2571 812
rect 2589 805 2594 812
rect 2711 805 2716 812
rect 2734 806 2739 813
rect 1831 656 1839 669
rect 2036 655 2042 660
rect 671 625 685 640
rect 2112 654 2117 659
rect 288 533 299 544
rect 2046 628 2051 633
rect 2122 627 2128 633
rect 2006 611 2012 617
rect 2133 616 2145 621
rect 2060 588 2065 593
rect 2214 611 2219 616
rect 2228 586 2233 591
rect 1459 547 1465 555
rect 1579 486 1585 493
rect 1539 472 1544 477
rect 1555 471 1560 476
rect 1571 471 1576 476
rect 2106 471 2111 476
rect 2038 446 2043 451
rect 1230 325 1239 331
rect 1271 389 1276 394
rect 1368 381 1373 386
rect 1418 388 1423 393
rect 1319 371 1326 378
rect 1514 379 1519 384
rect 1559 388 1564 393
rect 1360 356 1365 363
rect 1465 369 1472 376
rect 1650 379 1655 384
rect 1383 356 1388 363
rect 1278 345 1290 352
rect 1506 354 1511 361
rect 1529 354 1534 361
rect 1601 369 1608 376
rect 1642 354 1647 361
rect 1665 354 1670 361
rect 1439 335 1446 340
rect 1280 325 1289 332
rect 1642 335 1647 342
rect 1785 337 1792 344
rect 1727 328 1734 333
rect 1258 308 1271 316
rect 1439 295 1446 303
rect 1378 282 1383 287
rect 1276 239 1281 244
rect 1262 214 1267 219
rect 1229 193 1236 202
rect 1366 255 1372 261
rect 1343 244 1353 249
rect 1441 256 1446 261
rect 1430 216 1435 221
rect 1451 196 1458 202
rect 2115 444 2121 451
rect 1999 428 2004 433
rect 2129 433 2142 438
rect 2054 405 2059 410
rect 2208 428 2213 433
rect 2222 403 2227 408
rect 1716 282 1721 287
rect 1614 239 1619 244
rect 1600 214 1605 219
rect 1570 196 1577 202
rect 1706 255 1711 260
rect 1689 244 1700 249
rect 1779 256 1784 261
rect 1768 216 1773 221
rect 1366 179 1372 185
rect 1608 184 1615 190
rect 1706 180 1711 185
rect 1547 168 1554 176
rect 2094 299 2099 304
rect 2027 274 2032 279
rect 2102 272 2109 278
rect 1988 255 1993 261
rect 2115 261 2128 266
rect 2042 233 2047 238
rect 2196 256 2201 261
rect 2210 231 2215 236
rect 1547 -35 1553 -28
rect 1507 -49 1512 -44
rect 1523 -50 1528 -45
rect 1539 -50 1544 -45
rect 2085 115 2090 120
rect 2018 90 2023 95
rect 2094 88 2100 94
rect 1979 71 1984 78
rect 2106 77 2119 82
rect 2033 49 2038 54
rect 2187 72 2192 77
rect 2201 47 2206 52
rect 1198 -196 1207 -190
rect 1239 -132 1244 -127
rect 1336 -140 1341 -135
rect 1386 -133 1391 -128
rect 1287 -150 1294 -143
rect 1482 -142 1487 -137
rect 1527 -133 1532 -128
rect 1328 -165 1333 -158
rect 1433 -152 1440 -145
rect 1618 -142 1623 -137
rect 1351 -165 1356 -158
rect 1246 -176 1258 -169
rect 1474 -167 1479 -160
rect 1497 -167 1502 -160
rect 1569 -152 1576 -145
rect 1610 -167 1615 -160
rect 1633 -167 1638 -160
rect 1407 -186 1414 -181
rect 1248 -196 1257 -189
rect 1610 -186 1615 -179
rect 1753 -184 1760 -177
rect 1695 -193 1702 -188
rect 1226 -213 1239 -205
rect 1407 -226 1414 -218
rect 1346 -239 1351 -234
rect 1244 -282 1249 -277
rect 1230 -307 1235 -302
rect 1197 -328 1204 -319
rect 1334 -266 1340 -260
rect 1319 -277 1330 -272
rect 1409 -265 1414 -260
rect 1398 -305 1403 -300
rect 1419 -325 1426 -319
rect 1684 -239 1689 -234
rect 1582 -282 1587 -277
rect 1568 -307 1573 -302
rect 1538 -325 1545 -319
rect 1674 -266 1679 -261
rect 1657 -278 1669 -272
rect 1747 -265 1752 -260
rect 1736 -305 1741 -300
rect 1334 -342 1340 -336
rect 1576 -337 1583 -331
rect 1674 -341 1679 -336
rect 1515 -353 1522 -345
rect 1547 -486 1553 -479
rect 1507 -500 1512 -495
rect 1523 -501 1528 -496
rect 1539 -501 1544 -496
rect 1198 -647 1207 -641
rect 1239 -583 1244 -578
rect 1336 -591 1341 -586
rect 1386 -584 1391 -579
rect 1287 -601 1294 -594
rect 1482 -593 1487 -588
rect 1527 -584 1532 -579
rect 1328 -616 1333 -609
rect 1433 -603 1440 -596
rect 1618 -593 1623 -588
rect 1351 -616 1356 -609
rect 1246 -627 1258 -620
rect 1474 -618 1479 -611
rect 1497 -618 1502 -611
rect 1569 -603 1576 -596
rect 1610 -618 1615 -611
rect 1633 -618 1638 -611
rect 1407 -637 1414 -632
rect 1248 -647 1257 -640
rect 1610 -637 1615 -630
rect 1753 -635 1760 -628
rect 1695 -644 1702 -639
rect 1226 -664 1239 -656
rect 1407 -677 1414 -669
rect 1346 -690 1351 -685
rect 1244 -733 1249 -728
rect 1230 -758 1235 -753
rect 1197 -779 1204 -770
rect 1334 -717 1340 -711
rect 1319 -728 1330 -723
rect 1409 -716 1414 -711
rect 1398 -756 1403 -751
rect 1419 -776 1426 -770
rect 1684 -690 1689 -685
rect 1582 -733 1587 -728
rect 1568 -758 1573 -753
rect 1538 -776 1545 -770
rect 1674 -717 1679 -712
rect 1659 -728 1668 -723
rect 1747 -716 1752 -711
rect 1736 -756 1741 -751
rect 1334 -793 1340 -787
rect 1576 -788 1583 -782
rect 1674 -792 1679 -787
rect 1515 -804 1522 -796
rect 1554 -876 1565 -868
rect 1538 -936 1544 -929
rect 1498 -950 1503 -945
rect 1514 -951 1519 -946
rect 1530 -951 1535 -946
rect 1190 -1042 1200 -1032
rect 1189 -1097 1198 -1091
rect 1230 -1033 1235 -1028
rect 1327 -1041 1332 -1036
rect 1377 -1034 1382 -1029
rect 1278 -1051 1285 -1044
rect 1473 -1043 1478 -1038
rect 1518 -1034 1523 -1029
rect 1319 -1066 1324 -1059
rect 1424 -1053 1431 -1046
rect 1609 -1043 1614 -1038
rect 1342 -1066 1347 -1059
rect 1237 -1077 1249 -1070
rect 1465 -1068 1470 -1061
rect 1488 -1068 1493 -1061
rect 1560 -1053 1567 -1046
rect 1601 -1068 1606 -1061
rect 1624 -1068 1629 -1061
rect 1398 -1087 1405 -1082
rect 1239 -1097 1248 -1090
rect 1601 -1087 1606 -1080
rect 1744 -1085 1751 -1078
rect 1217 -1114 1230 -1106
rect 1398 -1127 1405 -1119
rect 1337 -1140 1342 -1135
rect 1235 -1183 1240 -1178
rect 1221 -1208 1226 -1203
rect 1188 -1229 1195 -1220
rect 1312 -1178 1321 -1173
rect 1400 -1166 1405 -1161
rect 1389 -1206 1394 -1201
rect 1410 -1226 1417 -1220
rect 1675 -1140 1680 -1135
rect 1573 -1183 1578 -1178
rect 1559 -1208 1564 -1203
rect 1529 -1226 1536 -1220
rect 1665 -1167 1670 -1162
rect 1648 -1178 1659 -1173
rect 1738 -1166 1743 -1161
rect 1727 -1206 1732 -1201
rect 1567 -1238 1574 -1232
rect 1665 -1242 1670 -1237
rect 1506 -1254 1513 -1246
<< metal2 >>
rect 918 1553 944 1556
rect 918 1549 923 1553
rect 902 1544 923 1549
rect 632 1528 936 1531
rect 632 1526 941 1528
rect 633 1447 636 1526
rect 869 1517 888 1522
rect 883 1469 888 1517
rect 944 1499 947 1517
rect 46 1444 636 1447
rect 46 1294 50 1444
rect 655 1426 669 1428
rect 872 1432 906 1437
rect 655 1424 674 1426
rect 707 1425 824 1428
rect 754 1424 824 1425
rect 655 1402 659 1424
rect 796 1402 800 1413
rect 342 1389 1071 1393
rect 125 1337 132 1342
rect 343 1321 348 1389
rect 554 1358 604 1362
rect 655 1362 660 1377
rect 742 1362 746 1389
rect 796 1364 800 1377
rect 931 1363 935 1379
rect 1925 1376 1932 1377
rect 1925 1375 2193 1376
rect 1925 1371 2194 1375
rect 571 1348 1257 1352
rect 199 1310 283 1318
rect 178 1302 234 1303
rect 86 1300 234 1302
rect 343 1300 349 1321
rect 86 1297 349 1300
rect 86 1296 184 1297
rect 45 1213 50 1294
rect 45 838 49 1213
rect 154 940 158 1273
rect 186 1049 189 1266
rect 229 1246 234 1297
rect 364 1294 461 1300
rect 364 1291 471 1294
rect 364 1271 369 1291
rect 361 1266 383 1271
rect 232 1223 250 1228
rect 288 1123 293 1240
rect 377 1228 383 1266
rect 390 1228 398 1233
rect 458 1228 463 1291
rect 571 1287 580 1348
rect 731 1331 840 1332
rect 645 1326 840 1331
rect 645 1325 759 1326
rect 538 1282 580 1287
rect 615 1312 655 1317
rect 681 1318 688 1325
rect 853 1326 856 1332
rect 1008 1327 1077 1330
rect 909 1325 1077 1327
rect 909 1322 1081 1325
rect 615 1281 621 1312
rect 796 1298 800 1315
rect 961 1283 966 1311
rect 1116 1264 1120 1325
rect 1177 1253 1182 1319
rect 1251 1307 1257 1348
rect 1925 1342 1932 1371
rect 1612 1336 1932 1342
rect 1955 1350 1960 1351
rect 1955 1344 2071 1350
rect 1177 1250 1206 1253
rect 556 1239 578 1245
rect 304 1158 309 1200
rect 462 1198 472 1202
rect 462 1158 468 1198
rect 556 1193 562 1239
rect 1177 1246 1185 1250
rect 1164 1241 1185 1246
rect 1250 1230 1257 1307
rect 1226 1227 1257 1230
rect 1226 1226 1254 1227
rect 1198 1221 1203 1225
rect 714 1199 720 1205
rect 561 1181 562 1193
rect 585 1180 739 1188
rect 304 1157 610 1158
rect 304 1153 612 1157
rect 633 1162 720 1163
rect 633 1156 721 1162
rect 457 1152 612 1153
rect 596 1150 612 1152
rect 517 1132 548 1139
rect 288 1118 570 1123
rect 186 892 189 1043
rect 226 1024 229 1072
rect 361 1069 468 1078
rect 361 1049 366 1069
rect 358 1044 380 1049
rect 229 1001 247 1006
rect 205 935 232 939
rect 161 888 189 892
rect 161 887 164 888
rect 152 881 164 887
rect 228 885 232 935
rect 287 916 291 1015
rect 374 1011 380 1044
rect 374 1006 379 1011
rect 455 1006 460 1069
rect 301 936 306 978
rect 459 976 469 980
rect 542 976 548 1091
rect 575 981 580 1064
rect 459 936 465 976
rect 301 933 465 936
rect 301 931 565 933
rect 454 930 565 931
rect 287 912 541 916
rect 398 897 480 901
rect 161 865 164 881
rect 200 882 232 885
rect 200 870 205 882
rect 186 867 205 870
rect 146 800 147 805
rect 146 782 149 800
rect 161 782 164 859
rect 186 805 190 867
rect 228 838 232 882
rect 364 884 471 893
rect 364 864 369 884
rect 361 859 383 864
rect 232 816 250 821
rect 161 778 189 782
rect 186 690 189 778
rect 228 663 231 788
rect 289 733 293 831
rect 377 821 383 859
rect 458 821 463 884
rect 304 751 309 793
rect 462 791 472 795
rect 462 751 468 791
rect 537 763 542 882
rect 560 861 565 930
rect 510 760 542 763
rect 510 759 541 760
rect 304 749 468 751
rect 558 750 565 861
rect 600 823 610 1150
rect 634 1124 640 1125
rect 634 1119 706 1124
rect 634 1021 640 1119
rect 699 1090 705 1119
rect 716 1106 721 1156
rect 758 1090 763 1205
rect 1613 1195 1621 1336
rect 1955 1322 1960 1344
rect 2188 1349 2194 1371
rect 2362 1364 3074 1368
rect 2371 1360 3074 1364
rect 802 1185 1621 1195
rect 781 1096 787 1112
rect 699 1086 763 1090
rect 780 1072 787 1096
rect 662 1065 787 1072
rect 620 1020 656 1021
rect 620 1019 664 1020
rect 620 1015 660 1019
rect 620 867 628 1015
rect 633 1014 660 1015
rect 733 1004 759 1007
rect 733 1000 738 1004
rect 717 995 738 1000
rect 803 984 810 1185
rect 1613 1184 1621 1185
rect 1635 1314 1960 1322
rect 1979 1318 2156 1323
rect 2188 1318 2193 1349
rect 2628 1327 2629 1336
rect 2246 1318 2456 1323
rect 1979 1317 2006 1318
rect 1635 1174 1641 1314
rect 943 1167 1642 1174
rect 815 1088 819 1110
rect 918 1088 923 1162
rect 815 1084 924 1088
rect 815 1019 819 1084
rect 880 1004 906 1007
rect 880 1000 885 1004
rect 864 995 885 1000
rect 779 981 810 984
rect 779 980 807 981
rect 751 961 756 979
rect 898 961 903 979
rect 943 983 950 1167
rect 1007 1156 1012 1162
rect 1024 1156 1039 1163
rect 959 1087 963 1093
rect 1007 1087 1014 1156
rect 1664 1145 1670 1295
rect 1980 1238 1986 1317
rect 2118 1310 2123 1311
rect 1892 1224 1918 1227
rect 1913 1220 1918 1224
rect 1913 1215 1934 1220
rect 1092 1140 1670 1145
rect 1772 1194 1777 1196
rect 1872 1195 1877 1199
rect 1855 1194 1877 1195
rect 1772 1190 1877 1194
rect 1772 1189 1861 1190
rect 1092 1137 1731 1140
rect 959 1081 1015 1087
rect 959 1017 963 1081
rect 1026 1002 1052 1005
rect 1026 998 1031 1002
rect 1010 993 1031 998
rect 926 979 950 983
rect 921 978 948 979
rect 1092 980 1097 1137
rect 1733 1136 1737 1137
rect 1253 1123 1260 1124
rect 1772 1123 1777 1189
rect 1253 1117 1777 1123
rect 1103 1096 1109 1101
rect 1103 1090 1199 1096
rect 1103 1014 1109 1090
rect 1162 1002 1188 1005
rect 1162 998 1167 1002
rect 1146 993 1167 998
rect 1072 977 1098 980
rect 1044 961 1049 977
rect 1180 961 1185 977
rect 1253 979 1260 1117
rect 1772 1115 1777 1117
rect 1208 977 1260 979
rect 1203 974 1260 977
rect 1318 1033 1323 1087
rect 1666 1056 1768 1060
rect 1585 1046 1611 1049
rect 1606 1042 1611 1046
rect 1606 1038 1627 1042
rect 1606 1037 1618 1038
rect 751 958 1270 961
rect 641 906 662 910
rect 724 897 750 900
rect 804 901 807 906
rect 724 893 729 897
rect 869 896 895 899
rect 708 888 729 893
rect 869 892 874 896
rect 853 887 874 892
rect 945 894 948 902
rect 1018 894 1044 897
rect 1018 890 1023 894
rect 1002 885 1023 890
rect 1090 883 1094 903
rect 1162 894 1188 897
rect 1162 890 1167 894
rect 1146 885 1167 890
rect 742 847 747 872
rect 770 872 792 876
rect 887 847 892 871
rect 915 871 931 873
rect 910 869 931 871
rect 1064 869 1074 873
rect 1036 847 1041 869
rect 1180 847 1185 869
rect 1208 868 1244 872
rect 1266 847 1270 958
rect 1318 904 1324 1033
rect 1433 1015 1488 1020
rect 1565 1020 1570 1022
rect 1496 1015 1570 1020
rect 1433 923 1438 1015
rect 1588 1005 1593 1023
rect 1520 998 1593 1005
rect 1433 921 1437 923
rect 1520 921 1527 998
rect 1584 928 1607 931
rect 1388 916 1405 921
rect 1435 916 1437 921
rect 1473 916 1527 921
rect 1602 924 1607 928
rect 1611 924 1616 1037
rect 1665 1037 1720 1043
rect 1671 937 1732 942
rect 1602 919 1624 924
rect 1318 897 1337 904
rect 1388 890 1394 916
rect 1442 899 1446 916
rect 1520 904 1527 916
rect 1520 903 1564 904
rect 1520 897 1569 903
rect 1586 890 1592 902
rect 1388 886 1592 890
rect 1388 885 1394 886
rect 742 844 1270 847
rect 742 843 747 844
rect 600 820 1090 823
rect 600 819 610 820
rect 896 799 900 804
rect 895 796 946 799
rect 953 796 954 799
rect 895 795 954 796
rect 772 781 805 784
rect 772 780 810 781
rect 558 749 616 750
rect 896 749 900 795
rect 1080 765 1247 771
rect 304 746 551 749
rect 289 729 502 733
rect 364 709 471 718
rect 510 709 516 715
rect 364 689 369 709
rect 361 684 383 689
rect 232 641 250 646
rect 288 561 292 656
rect 377 651 383 684
rect 377 646 378 651
rect 458 646 463 709
rect 304 576 309 618
rect 462 616 472 620
rect 462 577 468 616
rect 461 576 476 577
rect 304 571 476 576
rect 542 575 551 746
rect 558 746 903 749
rect 558 743 616 746
rect 940 749 1218 751
rect 940 745 1219 749
rect 800 717 1182 721
rect 626 628 671 637
rect 749 577 759 578
rect 631 576 759 577
rect 571 575 759 576
rect 542 572 759 575
rect 542 571 749 572
rect 1177 581 1182 717
rect 1209 614 1219 745
rect 1242 744 1247 765
rect 1242 666 1248 744
rect 1266 683 1270 844
rect 1319 710 1322 868
rect 1428 704 1432 886
rect 1583 824 1607 827
rect 1602 820 1607 824
rect 1611 820 1616 919
rect 1719 884 1722 937
rect 1763 902 1768 1056
rect 1792 1023 1795 1189
rect 1895 1183 1900 1199
rect 1991 1203 1996 1296
rect 2118 1239 2123 1303
rect 2151 1291 2156 1318
rect 2246 1291 2250 1318
rect 2028 1224 2054 1227
rect 2049 1220 2054 1224
rect 2049 1215 2070 1220
rect 1991 1199 2008 1203
rect 2134 1204 2139 1291
rect 2151 1287 2250 1291
rect 2264 1240 2269 1307
rect 2281 1288 2285 1292
rect 2281 1285 2402 1288
rect 2174 1226 2200 1229
rect 2195 1222 2200 1226
rect 2195 1217 2216 1222
rect 2134 1201 2154 1204
rect 2134 1200 2159 1201
rect 2139 1199 2155 1200
rect 1991 1198 2005 1199
rect 1991 1197 1996 1198
rect 2031 1183 2036 1199
rect 2177 1183 2182 1201
rect 2281 1206 2285 1285
rect 2421 1241 2427 1288
rect 2321 1226 2347 1229
rect 2342 1222 2347 1226
rect 2342 1217 2363 1222
rect 2289 1204 2297 1205
rect 2289 1201 2301 1204
rect 2289 1200 2306 1201
rect 2324 1183 2329 1201
rect 2450 1195 2456 1318
rect 2533 1225 2559 1228
rect 2554 1221 2559 1225
rect 2554 1216 2575 1221
rect 2513 1195 2518 1200
rect 2450 1190 2518 1195
rect 2625 1204 2629 1327
rect 2776 1304 2777 1313
rect 2669 1225 2695 1228
rect 2690 1221 2695 1225
rect 2690 1216 2711 1221
rect 2624 1200 2649 1204
rect 2771 1206 2777 1304
rect 2915 1286 2916 1293
rect 2815 1227 2841 1230
rect 2836 1223 2841 1227
rect 2836 1218 2857 1223
rect 2771 1205 2789 1206
rect 2771 1202 2795 1205
rect 2771 1201 2800 1202
rect 2911 1205 2916 1286
rect 2962 1227 2988 1230
rect 2983 1223 2988 1227
rect 2983 1218 3004 1223
rect 1810 1180 2329 1183
rect 1810 1069 1814 1180
rect 1892 1116 1918 1119
rect 1913 1112 1918 1116
rect 1993 1113 1998 1124
rect 2415 1127 2456 1132
rect 2036 1116 2062 1119
rect 1913 1107 1934 1112
rect 2057 1112 2062 1116
rect 2057 1107 2078 1112
rect 2133 1101 2139 1122
rect 2185 1118 2211 1121
rect 2206 1114 2211 1118
rect 2206 1109 2227 1114
rect 2284 1103 2288 1125
rect 2330 1119 2356 1122
rect 2351 1115 2356 1119
rect 2351 1110 2372 1115
rect 1861 1093 1872 1094
rect 1838 1090 1872 1093
rect 1895 1069 1900 1091
rect 2010 1091 2016 1094
rect 2010 1090 2021 1091
rect 2039 1069 2044 1091
rect 2159 1093 2165 1096
rect 2159 1092 2170 1093
rect 2188 1069 2193 1093
rect 2306 1093 2310 1097
rect 2333 1069 2338 1094
rect 1810 1066 2338 1069
rect 1810 1059 1814 1066
rect 2333 1065 2338 1066
rect 1806 1056 1814 1059
rect 1719 881 1772 884
rect 1669 833 1670 837
rect 1678 833 1719 837
rect 1602 815 1623 820
rect 1517 777 1545 782
rect 1583 728 1606 731
rect 1602 724 1606 728
rect 1611 726 1616 815
rect 1611 724 1612 726
rect 1602 719 1612 724
rect 1618 719 1624 724
rect 1428 701 1591 704
rect 1586 700 1591 701
rect 1713 683 1719 833
rect 1769 723 1772 881
rect 1806 743 1810 1056
rect 2154 1055 2158 1056
rect 1834 1028 1837 1051
rect 1833 847 1837 1028
rect 1848 1017 1854 1023
rect 2006 991 2010 1026
rect 2154 1001 2158 1049
rect 2364 1004 2367 1059
rect 2536 1023 2541 1200
rect 2672 1038 2677 1200
rect 2818 1054 2823 1202
rect 2910 1202 2942 1205
rect 2910 1201 2947 1202
rect 2965 1184 2970 1202
rect 2966 1135 2970 1184
rect 3067 1007 3074 1360
rect 1892 982 2010 991
rect 2153 992 2158 1001
rect 2177 999 2367 1004
rect 2528 1000 3074 1007
rect 1266 678 1719 683
rect 1713 677 1719 678
rect 1833 669 1837 841
rect 1892 817 1897 982
rect 1919 952 1928 954
rect 2153 952 2157 992
rect 1919 944 2160 952
rect 1243 638 1248 666
rect 1892 638 1897 809
rect 1919 759 1928 944
rect 2177 930 2189 999
rect 2369 947 2373 949
rect 2369 945 2377 947
rect 2373 942 2377 945
rect 2293 936 2319 939
rect 2314 932 2319 936
rect 1966 918 2189 930
rect 2223 927 2258 930
rect 2314 927 2335 932
rect 1926 751 1928 759
rect 1243 632 1902 638
rect 1209 609 1218 614
rect 1919 609 1928 751
rect 1967 724 1977 918
rect 2255 914 2258 927
rect 2255 911 2273 914
rect 2383 914 2386 993
rect 2511 945 2515 948
rect 2429 936 2455 939
rect 2450 932 2455 936
rect 2450 927 2471 932
rect 2383 911 2409 914
rect 2529 917 2534 1000
rect 2653 947 2655 951
rect 2825 946 2844 952
rect 2575 938 2601 941
rect 2596 934 2601 938
rect 2596 929 2617 934
rect 2529 913 2555 917
rect 2681 916 2685 940
rect 2722 938 2748 941
rect 2743 934 2748 938
rect 2743 929 2764 934
rect 2681 913 2702 916
rect 2296 895 2301 911
rect 2432 895 2437 911
rect 2578 895 2583 913
rect 2725 895 2730 913
rect 2211 892 2730 895
rect 2211 887 2215 892
rect 2104 884 2215 887
rect 2211 781 2215 884
rect 2372 837 2379 842
rect 2525 837 2534 841
rect 2674 839 2683 843
rect 2819 836 2822 845
rect 2293 828 2319 831
rect 2437 828 2463 831
rect 2586 830 2612 833
rect 2731 831 2757 834
rect 2314 824 2319 828
rect 2251 808 2254 824
rect 2314 819 2335 824
rect 2458 824 2463 828
rect 2607 826 2612 830
rect 2752 827 2757 831
rect 2458 819 2479 824
rect 2607 821 2628 826
rect 2752 822 2773 827
rect 2251 804 2273 808
rect 2296 781 2301 803
rect 2404 803 2417 807
rect 2422 803 2423 807
rect 2404 802 2423 803
rect 2552 805 2566 809
rect 2552 804 2571 805
rect 2690 806 2711 810
rect 2440 781 2445 803
rect 2589 781 2594 805
rect 2734 781 2739 806
rect 2211 778 2739 781
rect 2734 777 2739 778
rect 2007 761 2042 766
rect 1939 710 1943 717
rect 1209 599 1930 609
rect 1938 603 1943 710
rect 1919 597 1928 599
rect 1967 581 1977 716
rect 1177 572 1977 581
rect 2006 617 2010 689
rect 2036 660 2041 761
rect 2120 687 2227 688
rect 2120 684 2297 687
rect 2120 679 2227 684
rect 2120 659 2125 679
rect 2117 654 2139 659
rect 288 544 293 561
rect 1439 559 1466 564
rect 1459 555 1466 559
rect 1465 547 1466 555
rect 1579 493 1613 494
rect 1585 489 1613 493
rect 1273 473 1539 476
rect 1273 394 1276 473
rect 1555 467 1560 471
rect 1538 463 1560 467
rect 1538 452 1542 463
rect 1571 459 1576 471
rect 1419 447 1542 452
rect 1559 454 1576 459
rect 1419 393 1423 447
rect 1559 393 1563 454
rect 1342 381 1368 384
rect 1342 377 1347 381
rect 1326 372 1347 377
rect 1488 379 1514 382
rect 1619 382 1625 494
rect 1619 379 1650 382
rect 1488 375 1493 379
rect 1472 370 1493 375
rect 1619 375 1629 379
rect 1608 370 1629 375
rect 1210 345 1278 350
rect 1211 202 1215 345
rect 1239 325 1280 331
rect 1360 331 1365 356
rect 1383 339 1388 356
rect 1383 335 1439 339
rect 1506 339 1511 354
rect 1446 335 1511 339
rect 1529 339 1534 354
rect 1642 342 1647 354
rect 1529 335 1642 339
rect 1665 333 1670 354
rect 1727 333 1734 473
rect 1786 344 1792 474
rect 1882 465 1890 529
rect 2006 527 2011 611
rect 1884 428 1890 465
rect 1665 331 1727 333
rect 1360 328 1727 331
rect 1734 328 1784 333
rect 1271 308 1713 316
rect 1268 307 1713 308
rect 1276 244 1281 307
rect 1370 287 1375 307
rect 1356 282 1378 287
rect 1356 249 1362 282
rect 1441 261 1446 295
rect 1353 244 1362 249
rect 1267 214 1277 218
rect 1211 196 1229 202
rect 1271 174 1277 214
rect 1366 185 1372 255
rect 1614 244 1619 307
rect 1708 287 1713 307
rect 1694 282 1716 287
rect 1694 249 1700 282
rect 1779 261 1784 328
rect 1430 175 1435 216
rect 1605 214 1615 218
rect 1458 196 1570 202
rect 1609 190 1615 214
rect 1430 174 1547 175
rect 1271 170 1547 174
rect 1271 169 1435 170
rect 1609 174 1615 184
rect 1706 185 1711 255
rect 1768 174 1773 216
rect 1609 169 1773 174
rect 1882 138 1890 428
rect 1999 519 2011 527
rect 2046 603 2051 628
rect 2124 616 2128 627
rect 2133 621 2139 654
rect 2214 616 2219 679
rect 2120 613 2128 616
rect 2046 597 2047 603
rect 2046 526 2051 597
rect 2060 546 2065 588
rect 2218 586 2228 590
rect 2218 585 2232 586
rect 2218 549 2224 585
rect 2060 541 2216 546
rect 2293 532 2296 684
rect 2046 520 2050 526
rect 1999 433 2004 519
rect 2046 481 2051 520
rect 2293 513 2297 532
rect 1999 312 2004 428
rect 2038 478 2051 481
rect 2114 500 2221 505
rect 2293 500 2296 513
rect 2114 497 2297 500
rect 2114 496 2221 497
rect 2038 451 2043 478
rect 2114 476 2119 496
rect 2111 471 2133 476
rect 2038 364 2043 446
rect 2116 436 2120 444
rect 2127 438 2133 471
rect 2127 433 2129 438
rect 2208 433 2213 496
rect 1694 133 1890 138
rect 1988 308 2004 312
rect 2027 360 2043 364
rect 2054 363 2059 405
rect 2212 403 2222 407
rect 2212 402 2226 403
rect 2212 366 2218 402
rect 1988 261 1992 308
rect 2027 279 2032 360
rect 2054 358 2211 363
rect 2102 332 2209 333
rect 2293 332 2296 497
rect 2102 328 2296 332
rect 2102 324 2209 328
rect 2102 304 2107 324
rect 2099 299 2121 304
rect 1988 134 1992 255
rect 2027 188 2032 274
rect 2103 261 2107 272
rect 2115 266 2121 299
rect 2196 261 2201 324
rect 2018 185 2032 188
rect 2042 191 2047 233
rect 2200 231 2210 235
rect 2200 230 2214 231
rect 2200 193 2206 230
rect 2042 186 2199 191
rect 2018 144 2022 185
rect 2293 159 2296 328
rect 2291 150 2296 159
rect 2189 149 2296 150
rect 2093 145 2296 149
rect 1584 -27 1593 -26
rect 1547 -28 1593 -27
rect 1553 -32 1593 -28
rect 1584 -33 1593 -32
rect 1241 -48 1507 -45
rect 1241 -127 1244 -48
rect 1523 -54 1528 -50
rect 1506 -58 1528 -54
rect 1506 -69 1510 -58
rect 1539 -62 1544 -50
rect 1387 -74 1510 -69
rect 1527 -67 1544 -62
rect 1387 -128 1391 -74
rect 1527 -128 1531 -67
rect 1310 -140 1336 -137
rect 1310 -144 1315 -140
rect 1294 -149 1315 -144
rect 1456 -142 1482 -139
rect 1587 -139 1593 -33
rect 1587 -142 1618 -139
rect 1456 -146 1461 -142
rect 1440 -151 1461 -146
rect 1587 -146 1597 -142
rect 1576 -151 1597 -146
rect 1178 -176 1246 -171
rect 1179 -319 1183 -176
rect 1207 -196 1248 -190
rect 1328 -190 1333 -165
rect 1351 -182 1356 -165
rect 1351 -186 1407 -182
rect 1474 -182 1479 -167
rect 1414 -186 1479 -182
rect 1497 -182 1502 -167
rect 1610 -179 1615 -167
rect 1497 -186 1610 -182
rect 1633 -188 1638 -167
rect 1695 -188 1702 133
rect 1882 130 1890 133
rect 1979 130 1992 134
rect 2093 140 2200 145
rect 1979 78 1983 130
rect 2018 95 2022 133
rect 2093 120 2098 140
rect 2090 115 2112 120
rect 1978 71 1979 78
rect 2094 75 2098 88
rect 2106 82 2112 115
rect 2187 77 2192 140
rect 1978 70 1982 71
rect 2033 7 2038 49
rect 2191 47 2201 51
rect 2191 46 2205 47
rect 2191 9 2197 46
rect 2033 2 2191 7
rect 2186 1 2191 2
rect 1754 -53 1755 -44
rect 1767 -53 1772 -46
rect 1754 -177 1760 -53
rect 1633 -190 1695 -188
rect 1328 -193 1695 -190
rect 1702 -193 1752 -188
rect 1239 -213 1681 -205
rect 1236 -214 1681 -213
rect 1244 -277 1249 -214
rect 1338 -234 1343 -214
rect 1324 -239 1346 -234
rect 1324 -272 1330 -239
rect 1409 -260 1414 -226
rect 1235 -307 1245 -303
rect 1179 -325 1197 -319
rect 1239 -347 1245 -307
rect 1334 -336 1340 -266
rect 1582 -277 1587 -214
rect 1676 -234 1681 -214
rect 1662 -239 1684 -234
rect 1662 -272 1668 -239
rect 1747 -260 1752 -193
rect 1398 -346 1403 -305
rect 1573 -307 1583 -303
rect 1426 -325 1538 -319
rect 1577 -331 1583 -307
rect 1398 -347 1515 -346
rect 1239 -351 1515 -347
rect 1239 -352 1403 -351
rect 1577 -347 1583 -337
rect 1674 -336 1679 -266
rect 1736 -347 1741 -305
rect 1577 -352 1741 -347
rect 3103 -400 3116 985
rect 1695 -413 3117 -400
rect 1547 -479 1593 -478
rect 1553 -483 1593 -479
rect 1241 -499 1507 -496
rect 1241 -578 1244 -499
rect 1523 -505 1528 -501
rect 1506 -509 1528 -505
rect 1506 -520 1510 -509
rect 1539 -513 1544 -501
rect 1387 -525 1510 -520
rect 1527 -518 1544 -513
rect 1387 -579 1391 -525
rect 1527 -579 1531 -518
rect 1310 -591 1336 -588
rect 1310 -595 1315 -591
rect 1294 -600 1315 -595
rect 1456 -593 1482 -590
rect 1587 -590 1593 -483
rect 1696 -494 1702 -413
rect 1587 -593 1618 -590
rect 1456 -597 1461 -593
rect 1440 -602 1461 -597
rect 1587 -597 1597 -593
rect 1576 -602 1597 -597
rect 1178 -627 1246 -622
rect 1179 -770 1183 -627
rect 1207 -647 1248 -641
rect 1328 -641 1333 -616
rect 1351 -633 1356 -616
rect 1351 -637 1407 -633
rect 1474 -633 1479 -618
rect 1414 -637 1479 -633
rect 1497 -633 1502 -618
rect 1610 -630 1615 -618
rect 1497 -637 1610 -633
rect 1633 -639 1638 -618
rect 1695 -639 1702 -494
rect 1754 -628 1760 -499
rect 1850 -552 1928 -542
rect 1633 -641 1695 -639
rect 1328 -644 1695 -641
rect 1702 -644 1752 -639
rect 1239 -664 1681 -656
rect 1236 -665 1681 -664
rect 1244 -728 1249 -665
rect 1338 -685 1343 -665
rect 1324 -690 1346 -685
rect 1324 -723 1330 -690
rect 1409 -711 1414 -677
rect 1235 -758 1245 -754
rect 1179 -776 1197 -770
rect 1239 -798 1245 -758
rect 1334 -787 1340 -717
rect 1582 -728 1587 -665
rect 1676 -685 1681 -665
rect 1662 -690 1684 -685
rect 1662 -723 1668 -690
rect 1747 -711 1752 -644
rect 1398 -797 1403 -756
rect 1573 -758 1583 -754
rect 1426 -776 1538 -770
rect 1577 -782 1583 -758
rect 1398 -798 1515 -797
rect 1239 -802 1515 -798
rect 1239 -803 1403 -802
rect 1577 -798 1583 -788
rect 1674 -787 1679 -717
rect 1736 -798 1741 -756
rect 1577 -803 1741 -798
rect 1194 -830 1200 -829
rect 1850 -830 1857 -552
rect 1194 -836 1857 -830
rect 1194 -1032 1200 -836
rect 1589 -870 1607 -869
rect 1565 -876 1607 -870
rect 1589 -877 1607 -876
rect 1618 -877 1620 -869
rect 3209 -911 3221 1048
rect 1686 -918 3224 -911
rect 1538 -929 1584 -928
rect 1544 -933 1584 -929
rect 1232 -949 1498 -946
rect 1232 -1028 1235 -949
rect 1514 -955 1519 -951
rect 1497 -959 1519 -955
rect 1497 -970 1501 -959
rect 1530 -963 1535 -951
rect 1378 -975 1501 -970
rect 1518 -968 1535 -963
rect 1378 -1029 1382 -975
rect 1518 -1029 1522 -968
rect 1301 -1041 1327 -1038
rect 1301 -1045 1306 -1041
rect 1285 -1050 1306 -1045
rect 1447 -1043 1473 -1040
rect 1578 -1040 1584 -933
rect 1687 -944 1695 -918
rect 1686 -960 1695 -944
rect 1578 -1043 1609 -1040
rect 1447 -1047 1452 -1043
rect 1431 -1052 1452 -1047
rect 1578 -1047 1588 -1043
rect 1567 -1052 1588 -1047
rect 1169 -1077 1237 -1072
rect 1170 -1220 1174 -1077
rect 1198 -1097 1239 -1091
rect 1319 -1091 1324 -1066
rect 1342 -1083 1347 -1066
rect 1342 -1087 1398 -1083
rect 1465 -1083 1470 -1068
rect 1405 -1087 1470 -1083
rect 1488 -1083 1493 -1068
rect 1601 -1080 1606 -1068
rect 1488 -1087 1601 -1083
rect 1624 -1089 1629 -1068
rect 1686 -1089 1693 -960
rect 1745 -1078 1751 -946
rect 1624 -1091 1743 -1089
rect 1319 -1094 1743 -1091
rect 1230 -1114 1672 -1106
rect 1219 -1115 1672 -1114
rect 1235 -1178 1240 -1115
rect 1329 -1135 1334 -1115
rect 1315 -1140 1337 -1135
rect 1315 -1173 1321 -1140
rect 1400 -1161 1405 -1127
rect 1573 -1178 1578 -1115
rect 1667 -1135 1672 -1115
rect 1653 -1140 1675 -1135
rect 1653 -1173 1659 -1140
rect 1738 -1161 1743 -1094
rect 1226 -1208 1236 -1204
rect 1170 -1226 1188 -1220
rect 1230 -1248 1236 -1208
rect 1389 -1247 1394 -1206
rect 1564 -1208 1574 -1204
rect 1417 -1226 1529 -1220
rect 1568 -1232 1574 -1208
rect 1389 -1248 1506 -1247
rect 1230 -1252 1506 -1248
rect 1230 -1253 1394 -1252
rect 1568 -1248 1574 -1238
rect 1665 -1237 1670 -1167
rect 1727 -1248 1732 -1206
rect 1568 -1253 1732 -1248
<< m3contact >>
rect 906 1431 913 1437
rect 824 1421 837 1429
rect 113 1334 125 1346
rect 546 1357 554 1366
rect 283 1309 299 1321
rect 152 1273 160 1281
rect 631 1323 645 1334
rect 1114 1325 1127 1332
rect 959 1311 967 1316
rect 1197 1215 1205 1221
rect 706 1199 714 1207
rect 387 897 398 905
rect 1731 1137 1737 1142
rect 1199 1090 1207 1096
rect 804 896 809 901
rect 945 889 950 894
rect 1090 878 1095 883
rect 792 872 797 878
rect 931 868 938 874
rect 1074 869 1080 876
rect 1090 819 1095 824
rect 946 796 953 802
rect 763 779 772 787
rect 805 781 812 787
rect 1072 765 1080 775
rect 510 715 517 723
rect 931 745 940 754
rect 795 717 800 725
rect 759 569 771 582
rect 2402 1285 2407 1291
rect 2421 1288 2429 1296
rect 2906 1286 2915 1296
rect 2456 1125 2466 1133
rect 1993 1107 1998 1113
rect 2004 1088 2010 1096
rect 2132 1094 2139 1101
rect 2153 1089 2159 1097
rect 2283 1096 2289 1103
rect 2298 1091 2306 1101
rect 2361 1059 2368 1065
rect 1507 773 1517 784
rect 1612 719 1618 726
rect 2153 1049 2160 1055
rect 1848 1023 1855 1030
rect 2004 1026 2012 1033
rect 2965 1126 2975 1135
rect 2816 1046 2826 1054
rect 2669 1031 2679 1038
rect 2536 1015 2543 1023
rect 3207 1048 3231 1069
rect 1833 841 1839 847
rect 1891 809 1898 817
rect 2373 937 2378 942
rect 1917 751 1926 759
rect 2515 944 2520 949
rect 3100 985 3122 1002
rect 2655 946 2661 951
rect 2681 940 2686 945
rect 2844 944 2851 954
rect 2379 837 2385 842
rect 2534 837 2539 842
rect 2683 839 2688 844
rect 2251 824 2256 829
rect 2817 831 2822 836
rect 2397 802 2404 807
rect 2547 804 2552 809
rect 2684 806 2690 811
rect 1966 716 1977 724
rect 1938 597 1945 603
rect 1430 558 1439 566
rect 1875 529 1896 537
rect 1613 488 1619 495
rect 1725 473 1738 483
rect 1786 474 1797 483
rect 2114 613 2120 618
rect 2047 597 2053 603
rect 2216 541 2224 549
rect 2116 431 2121 436
rect 2211 358 2218 366
rect 2102 256 2109 261
rect 2199 185 2207 193
rect 2014 133 2025 144
rect 2093 70 2099 75
rect 2191 1 2199 9
rect 1755 -53 1767 -42
rect 1754 -499 1766 -482
rect 1928 -560 1941 -538
rect 1607 -878 1618 -869
rect 1744 -946 1758 -934
<< metal3 >>
rect 913 1431 1033 1436
rect 1029 1422 1033 1431
rect 829 1419 1000 1421
rect 1029 1419 1119 1422
rect 829 1417 1001 1419
rect 1029 1417 1121 1419
rect 154 1364 157 1365
rect 152 1359 546 1364
rect 116 926 120 1334
rect 154 1281 157 1359
rect 390 1330 394 1332
rect 535 1330 631 1331
rect 389 1326 631 1330
rect 390 1318 394 1326
rect 535 1324 631 1326
rect 299 1309 395 1318
rect 997 1316 1001 1417
rect 1116 1332 1121 1417
rect 2402 1374 3087 1378
rect 967 1311 1002 1316
rect 2402 1291 2406 1374
rect 2429 1294 2439 1295
rect 2429 1289 2906 1294
rect 2429 1288 2439 1289
rect 607 1134 615 1136
rect 707 1134 712 1199
rect 606 1127 713 1134
rect 580 943 587 945
rect 607 943 615 1127
rect 1199 1096 1202 1215
rect 1733 1096 1737 1137
rect 2461 1133 2965 1135
rect 2466 1126 2965 1133
rect 1781 1100 1852 1103
rect 1781 1096 1785 1100
rect 1733 1092 1785 1096
rect 1848 1030 1852 1100
rect 1993 1018 1998 1107
rect 2005 1033 2010 1088
rect 2132 1038 2139 1094
rect 2154 1055 2158 1089
rect 2283 1051 2289 1096
rect 2300 1063 2303 1091
rect 2300 1060 2361 1063
rect 2283 1046 2816 1051
rect 2132 1032 2669 1038
rect 1993 1015 2536 1018
rect 3081 1019 3087 1374
rect 3139 1048 3207 1060
rect 2673 1015 3087 1019
rect 1993 1014 2542 1015
rect 2661 946 2664 951
rect 580 936 616 943
rect 2378 937 2380 940
rect 116 922 248 926
rect 240 902 245 922
rect 240 898 387 902
rect 580 825 587 936
rect 1725 922 1732 925
rect 1725 917 2265 922
rect 797 872 798 877
rect 579 721 587 825
rect 517 715 587 721
rect 761 779 763 785
rect 761 582 766 779
rect 795 725 798 872
rect 806 787 809 896
rect 931 754 937 868
rect 946 802 949 889
rect 1073 869 1074 871
rect 1073 775 1079 869
rect 1090 824 1094 878
rect 1430 780 1507 781
rect 1429 776 1507 780
rect 1101 567 1203 568
rect 1429 567 1436 776
rect 1517 776 1518 781
rect 1098 566 1203 567
rect 1400 566 1436 567
rect 1098 565 1271 566
rect 1400 565 1430 566
rect 1098 560 1430 565
rect 1098 165 1108 560
rect 1169 558 1430 560
rect 1233 557 1416 558
rect 1613 495 1618 719
rect 1725 483 1732 917
rect 2262 907 2265 917
rect 2376 907 2380 937
rect 2515 939 2519 944
rect 2659 937 2664 946
rect 2673 945 2676 1015
rect 3085 999 3100 1001
rect 3078 985 3100 999
rect 3078 984 3107 985
rect 2844 954 2851 971
rect 2673 941 2681 945
rect 3078 961 3089 984
rect 3063 950 3089 961
rect 2659 934 2666 937
rect 2262 903 2380 907
rect 1839 841 2254 845
rect 2251 829 2254 841
rect 2381 829 2385 837
rect 2534 827 2538 837
rect 2684 831 2688 839
rect 2819 822 2822 831
rect 1898 809 2188 814
rect 1880 793 1890 800
rect 1884 537 1889 793
rect 2182 770 2188 809
rect 2399 770 2404 802
rect 2182 764 2404 770
rect 2547 757 2552 804
rect 1926 751 2552 757
rect 2684 724 2689 806
rect 1977 716 2689 724
rect 1945 597 2047 603
rect 1786 518 1792 519
rect 2114 518 2118 613
rect 2224 541 2379 546
rect 1786 512 2119 518
rect 1786 483 1792 512
rect 2121 431 2122 435
rect 2119 342 2122 431
rect 2218 358 2402 363
rect 1858 337 2122 342
rect 1096 119 1108 165
rect 1096 -165 1106 119
rect 1859 -46 1869 337
rect 2103 164 2108 256
rect 2207 187 2418 192
rect 1767 -53 1869 -46
rect 1907 157 2108 164
rect 1094 -283 1106 -165
rect 1094 -836 1104 -283
rect 1907 -484 1916 157
rect 1766 -494 1916 -484
rect 1930 133 2014 142
rect 1930 -538 1937 133
rect 2093 75 2097 78
rect 1094 -846 1550 -836
rect 1094 -851 1618 -846
rect 1541 -853 1618 -851
rect 1610 -869 1618 -853
rect 2093 -938 2097 70
rect 2378 6 2384 7
rect 2199 2 2444 6
rect 1861 -939 2097 -938
rect 1758 -946 2097 -939
rect 2093 -947 2097 -946
<< m4contact >>
rect 3122 1048 3139 1067
rect 2515 934 2520 939
rect 2842 971 2853 980
rect 3047 950 3063 970
rect 2666 931 2674 937
rect 2381 824 2386 829
rect 2534 822 2539 827
rect 2683 826 2689 831
rect 2818 817 2823 822
rect 1871 792 1880 803
rect 2379 541 2384 546
rect 2402 358 2408 365
rect 2418 186 2426 193
rect 2444 0 2450 8
<< metal4 >>
rect 2845 1083 2852 1084
rect 2845 1075 2953 1083
rect 2845 980 2852 1075
rect 2945 1063 2953 1075
rect 2945 1052 3122 1063
rect 2874 959 2882 960
rect 2872 950 3047 959
rect 2872 949 3062 950
rect 2874 944 2882 949
rect 2505 934 2515 937
rect 2505 900 2508 934
rect 2195 895 2509 900
rect 2668 899 2672 931
rect 2874 909 2883 944
rect 2875 900 2883 909
rect 2785 899 2884 900
rect 2195 825 2199 895
rect 2668 891 2884 899
rect 2668 890 2807 891
rect 2381 829 2385 836
rect 1870 820 2201 825
rect 1871 803 1881 820
rect 2195 819 2199 820
rect 1880 792 1881 803
rect 2381 546 2385 824
rect 2685 822 2689 826
rect 2384 541 2385 546
rect 2381 533 2385 541
rect 2380 526 2385 533
rect 2402 695 2407 696
rect 2534 695 2538 822
rect 2685 819 2699 822
rect 2694 704 2699 819
rect 2820 778 2823 817
rect 2750 777 2823 778
rect 2749 774 2823 777
rect 2749 766 2753 774
rect 2820 773 2823 774
rect 2402 691 2538 695
rect 2549 699 2699 704
rect 2707 762 2754 766
rect 2402 526 2407 691
rect 2549 677 2554 699
rect 2707 685 2710 762
rect 2419 673 2554 677
rect 2572 681 2710 685
rect 2419 672 2553 673
rect 2419 526 2424 672
rect 2572 659 2575 681
rect 2445 655 2575 659
rect 2380 520 2384 526
rect 2402 520 2406 526
rect 2419 520 2423 526
rect 2380 514 2385 520
rect 2381 -5 2385 514
rect 2402 442 2407 520
rect 2401 365 2407 442
rect 2401 358 2402 365
rect 2401 60 2406 358
rect 2419 193 2424 520
rect 2419 137 2424 186
rect 2401 29 2407 60
rect 2402 -5 2407 29
rect 2418 56 2424 137
rect 2418 -5 2423 56
rect 2445 8 2449 655
<< labels >>
rlabel metal1 1426 919 1426 919 1 S0c
rlabel metal1 1411 919 1411 919 1 S0
rlabel metal1 1449 920 1449 920 1 S1
rlabel metal1 1665 939 1665 939 1 D1
rlabel metal1 1659 1058 1659 1058 1 D0
rlabel metal1 1667 739 1667 739 1 D3
rlabel metal1 1576 722 1576 722 1 DEC_AND_NODE_4
rlabel metal1 1576 745 1576 745 1 DEC_D3_NAND
rlabel metal1 1668 835 1668 835 1 D2
rlabel metal1 1577 818 1577 818 1 DEC_AND_NODE_3
rlabel metal1 1577 841 1577 841 1 DEC_D2_NAND
rlabel metal1 1579 922 1579 922 1 Dec_AND_node_2
rlabel metal1 1580 945 1580 945 1 DEC_D1_NAND
rlabel metal1 1575 1064 1575 1064 1 DEC_D0_NAND
rlabel metal1 1580 1041 1580 1041 1 Dec_AND_node_1
rlabel m2contact 1468 919 1468 919 1 S1c
rlabel metal1 1468 901 1468 901 1 gnd
rlabel metal1 1444 945 1444 945 1 vdd
rlabel metal2 1867 1092 1867 1092 1 B3
rlabel m3contact 2008 1093 2008 1093 1 B2
rlabel metal2 2160 1095 2160 1095 1 B1
rlabel metal1 2326 1113 2326 1113 1 ander_node_5
rlabel metal1 2178 1113 2178 1113 1 ander_node_6
rlabel metal1 2029 1109 2029 1109 1 ander_node_7
rlabel metal1 1884 1111 1884 1111 1 ander_node_8
rlabel metal1 2360 1130 2360 1130 1 and_b0e_nand
rlabel metal1 2225 1129 2225 1129 1 and_b1e_nand
rlabel metal1 2071 1126 2071 1126 1 and_b2e_nand
rlabel metal1 1923 1126 1923 1126 1 and_b3e_nand
rlabel metal1 2404 1130 2404 1130 1 and_b0e
rlabel metal1 2260 1129 2260 1129 1 and_b1e
rlabel metal1 2112 1126 2112 1126 1 and_b2e
rlabel metal1 1968 1127 1968 1127 1 and_b3e
rlabel metal1 2395 1236 2395 1236 1 and_a0e
rlabel metal1 2248 1236 2248 1236 1 and_a1e
rlabel metal1 2101 1234 2101 1234 1 and_a2e
rlabel metal1 1966 1235 1966 1235 1 and_a3e
rlabel metal1 2358 1236 2358 1236 1 and_a0e_nand
rlabel metal1 2212 1237 2212 1237 1 and_a1e_nand
rlabel metal1 2069 1235 2069 1235 1 and_a2e_nand
rlabel metal1 1925 1236 1925 1236 1 and_a3e_nand
rlabel metal1 2315 1220 2315 1220 1 ander_node_4
rlabel metal1 2168 1220 2168 1220 1 ander_node_3
rlabel metal1 2022 1219 2022 1219 1 ander_node_2
rlabel metal1 1886 1218 1886 1218 1 ander_node_1
rlabel metal2 2295 1202 2295 1202 1 A0
rlabel metal2 2149 1202 2149 1202 1 A1
rlabel metal2 2002 1200 2002 1200 1 A2
rlabel metal2 1874 1195 1874 1195 1 A3
rlabel metal1 2526 1220 2526 1220 1 ander_node_9
rlabel metal1 2660 1220 2660 1220 1 ander_node_10
rlabel metal1 2810 1223 2810 1223 1 ander_node_11
rlabel metal1 2954 1220 2954 1220 1 ander_node_12
rlabel metal1 2567 1236 2567 1236 1 A3_and_B3_nand
rlabel metal1 2695 1237 2695 1237 1 A2_and_B2_nand
rlabel metal1 2850 1238 2850 1238 1 A1_and_B1_nand
rlabel metal1 2990 1238 2990 1238 1 A0_and_B0_nand
rlabel metal1 2608 1236 2608 1236 1 A3_and_B3
rlabel metal1 2744 1236 2744 1236 1 A2_and_B2
rlabel metal1 2889 1238 2889 1238 1 A1_and_B1
rlabel metal1 3037 1238 3037 1238 1 A0_and_B0
rlabel metal1 1197 997 1197 997 1 compare_node_1
rlabel metal1 1058 997 1058 997 1 compare_node_2
rlabel metal1 912 998 912 998 1 compare_node_3
rlabel metal1 766 998 766 998 1 compare_node_4
rlabel metal1 757 892 757 892 1 compare_node_5
rlabel metal1 901 890 901 890 1 compare_node_6
rlabel metal1 1051 887 1051 887 1 compare_node_7
rlabel metal1 1194 887 1194 887 1 compare_node_8
rlabel metal1 1197 1028 1197 1028 1 compare_A3e_nand
rlabel metal1 1063 1027 1063 1027 1 compare_A2e_nand
rlabel metal1 917 1026 917 1026 1 compare_A1e_nand
rlabel metal1 769 1030 769 1030 1 compare_A0e_nand
rlabel metal1 761 923 761 923 1 compare_B0e_nand
rlabel metal1 906 920 906 920 1 compare_B1e_nand
rlabel metal1 1054 919 1054 919 1 compare_B2e_nand
rlabel metal1 1199 919 1199 919 1 compare_B3e_nand
rlabel metal1 1113 1013 1113 1013 1 compare_A3e
rlabel metal1 978 1014 978 1014 1 compare_A2e
rlabel metal1 834 1014 834 1014 1 compare_A1e
rlabel metal1 685 1016 685 1016 1 compare_A0e
rlabel metal1 677 908 677 908 1 compare_B0e
rlabel metal1 823 907 823 907 1 compare_B1e
rlabel metal1 972 904 972 904 1 compare_B2e
rlabel metal1 1117 905 1117 905 1 compare_B3e
rlabel pdiffusion 335 1253 335 1253 1 xnor_1
rlabel ndiffusion 335 1213 335 1213 1 xnor_2
rlabel metal1 396 1242 396 1242 1 xor_1
rlabel ndiffusion 417 1253 417 1253 1 xnor_3
rlabel pdiffusion 417 1213 417 1213 1 xnor_4
rlabel metal1 425 1167 425 1167 1 A3c
rlabel metal1 382 1284 382 1284 1 B3c
rlabel pdiffusion 330 1031 330 1031 1 xnor_5
rlabel ndiffusion 333 991 333 991 1 xnor_6
rlabel ndiffusion 416 1031 416 1031 1 xnor_7
rlabel pdiffusion 412 990 412 990 1 xnor_8
rlabel metal1 424 942 424 942 1 A2c
rlabel metal1 383 1064 383 1064 1 B2c
rlabel metal1 383 879 383 879 1 B1c
rlabel metal1 417 756 417 756 1 A1c
rlabel pdiffusion 335 845 335 845 1 xnor_9
rlabel ndiffusion 338 806 338 806 1 xnor_10
rlabel pdiffusion 416 806 416 806 1 xnor_11
rlabel ndiffusion 418 846 418 846 1 xnor_12
rlabel metal1 385 1018 385 1018 1 xor_2
rlabel metal1 390 834 390 834 1 xor_3
rlabel metal1 393 703 393 703 1 B0c
rlabel metal1 417 582 417 582 1 A0c
rlabel metal1 393 660 393 660 1 xor_4
rlabel pdiffusion 334 671 334 671 1 xnor_13
rlabel ndiffusion 336 630 336 630 1 xnor_14
rlabel ndiffusion 418 670 418 670 1 xnor_15
rlabel pdiffusion 418 631 418 631 1 xnor_16
rlabel ndiffusion 88 823 88 823 1 A_compare_B_node_3
rlabel ndiffusion 105 824 105 824 1 A_compare_B_node_2
rlabel ndiffusion 120 824 120 824 1 A_compare_B_node_1
rlabel metal1 5 848 5 848 3 A_equal_B
rlabel metal1 51 836 51 836 1 A_equal_B_c
rlabel metal1 94 906 94 906 1 A2e_xnor_B2e
rlabel metal1 223 1244 223 1244 1 A3e_xnor_B3e
rlabel metal1 222 836 222 836 1 A1e_xnor_B1e
rlabel metal1 223 660 223 660 1 A0e_xnor_B0e
rlabel metal2 2307 1094 2307 1094 1 B0
rlabel metal1 1214 1245 1214 1245 1 A_greater_B_node_1
rlabel metal1 1126 1261 1126 1261 1 A3_and_B3c
rlabel metal1 1211 1277 1211 1277 1 A3_nand_B3c
rlabel ndiffusion 1070 1253 1070 1253 1 A_greater_B_node_2
rlabel ndiffusion 1054 1253 1054 1253 1 A_greater_B_node_3
rlabel metal1 1024 1261 1024 1261 1 A3_eq_B3_A2_gt_B2_c
rlabel metal1 969 1279 969 1279 1 A3_eq_B3_A2_gt_B2
rlabel ndiffusion 928 1254 928 1254 1 A_greater_B_node_5
rlabel ndiffusion 907 1255 907 1255 1 A_greater_B_node_6
rlabel ndiffusion 891 1253 891 1253 1 A_greater_B_node_7
rlabel metal1 866 1267 866 1267 1 A3_eq_B3_A2_eq_B2_A1_gt_B1_c
rlabel metal1 812 1280 812 1280 1 A3_eq_B3_A2_eq_B2_A1_gt_B1
rlabel ndiffusion 734 1256 734 1256 1 A_greater_B_node_9
rlabel ndiffusion 715 1255 715 1255 1 A_greater_B_node_10
rlabel ndiffusion 699 1255 699 1255 1 A_greater_B_node_11
rlabel metal1 675 1265 675 1265 1 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c
rlabel metal1 622 1279 622 1279 1 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0
rlabel ndiffusion 750 1254 750 1254 1 A_greater_B_node_8
rlabel pdiffusion 710 1492 710 1492 1 A_GT_B_node_1
rlabel pdiffusion 694 1491 694 1491 1 A_GT_B_node_2
rlabel pdiffusion 677 1493 677 1493 1 A_GT_B_node_3
rlabel metal1 750 1466 750 1466 1 A_GT_B_c
rlabel metal1 792 1483 792 1483 1 A_GT_B
rlabel metal1 948 1547 948 1547 1 A_LS_B_node_1
rlabel metal1 954 1578 954 1578 1 A_LS_B_nand
rlabel metal1 864 1564 864 1564 1 A_LS_B
rlabel metal1 2028 872 2028 872 1 D0_OR_D1_node
rlabel metal1 2027 898 2027 898 1 D0_OR_D1_node_2
rlabel metal1 2063 882 2063 882 1 D0_or_D1_c
rlabel metal1 2096 886 2096 886 1 D0_or_D1
rlabel metal1 2286 930 2286 930 1 adder_node1
rlabel metal1 2421 931 2421 931 1 adder_node2
rlabel metal1 2565 933 2565 933 1 adder_node3
rlabel metal1 2716 932 2716 932 1 adder_node4
rlabel metal1 2724 825 2724 825 1 adder_node5
rlabel metal1 2585 823 2585 823 1 adder_node6
rlabel metal1 2430 823 2430 823 1 adder_node7
rlabel metal1 2285 821 2285 821 1 adder_node8
rlabel metal1 2324 947 2324 947 1 Adder_A3ec
rlabel metal1 2463 946 2463 946 1 Adder_A2ec
rlabel metal1 2619 949 2619 949 1 Adder_A1ec
rlabel metal1 2754 948 2754 948 1 Adder_A0ec
rlabel metal1 2763 841 2763 841 1 Adder_B0ec
rlabel metal1 2635 840 2635 840 1 Adder_B1ec
rlabel metal1 2474 839 2474 839 1 Adder_B2ec
rlabel metal1 2325 839 2325 839 1 Adder_B3ec
rlabel metal1 2366 947 2366 947 1 adder_A3e
rlabel metal1 2502 946 2502 946 1 adder_A2e
rlabel metal1 2648 948 2648 948 1 adder_A1e
rlabel metal1 2795 948 2795 948 1 adder_A0e
rlabel metal1 2803 841 2803 841 1 adder_B0e
rlabel metal1 2661 840 2661 840 1 adder_B1e
rlabel metal1 2511 838 2511 838 1 adder_B2e
rlabel metal1 2367 839 2367 839 1 adder_B3e
rlabel metal1 2186 673 2186 673 1 B3ec_M
rlabel metal1 2186 490 2186 490 1 B2ec_M
rlabel metal1 2217 317 2217 317 1 B1ec_M
rlabel metal1 2235 135 2235 135 1 01ec_M
rlabel ndiffusion 2171 640 2171 640 1 adder_xor_node1
rlabel pdiffusion 2089 641 2089 641 1 adder_xor_node2
rlabel pdiffusion 2175 602 2175 602 1 adder_xor_node4
rlabel pdiffusion 2085 458 2085 458 1 adder_xor_node5
rlabel ndiffusion 2167 458 2167 458 1 adder_xor_node6
rlabel ndiffusion 2082 420 2082 420 1 adder_xor_node7
rlabel pdiffusion 2166 419 2166 419 1 adder_xor_node8
rlabel ndiffusion 2155 284 2155 284 1 adder_xor_node9
rlabel pdiffusion 2071 284 2071 284 1 adder_xor_node10
rlabel ndiffusion 2073 248 2073 248 1 adder_xor_node11
rlabel pdiffusion 2159 245 2159 245 1 adder_xor_node12
rlabel pdiffusion 2062 101 2062 101 1 adder_xor_node13
rlabel ndiffusion 2145 102 2145 102 1 adder_xor_node14
rlabel ndiffusion 2063 62 2063 62 1 adder_xor_node15
rlabel pdiffusion 2146 61 2146 61 1 adder_xor_node16
rlabel metal1 2119 629 2119 629 1 B3e_xor_M
rlabel metal1 2103 434 2103 434 1 B2e_xor_M
rlabel metal1 2090 266 2090 266 1 B1e_xor_M
rlabel metal1 2079 79 2079 79 1 B0e_xor_M
rlabel ndiffusion 2093 601 2093 601 1 adder_xor_node3
rlabel metal1 1402 -897 1402 -897 1 carry1
rlabel metal2 1337 -741 1337 -741 1 Sum1
rlabel metal1 1389 -448 1389 -448 1 carry2
rlabel metal2 1336 -300 1336 -300 1 sum2
rlabel metal1 1377 3 1377 3 1 carry3
rlabel metal2 1367 235 1367 235 1 sum3
rlabel metal1 1430 526 1430 526 1 sum4
rlabel metal1 1329 -1163 1329 -1163 1 Sum0
rlabel metal1 1647 -1166 1647 -1166 1 A0_B0_XOR
<< end >>
