* SPICE3 file created from DECODER.ext - technology: scmos

.option scale=90n

M1000 DEC_D1_NAND S1c vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1001 vdd S0 DEC_D1_NAND vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1002 DEC_D2_NAND S0c DEC_AND_NODE_3 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1003 Dec_AND_node_1 S1c gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1004 DEC_AND_NODE_3 S1 gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1005 S1c S1 vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1006 S0c S0 gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1007 D0 DEC_D0_NAND gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1008 DEC_D3_NAND S1 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1009 D3 DEC_D3_NAND vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1010 DEC_D1_NAND S1c Dec_AND_node_2 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1011 Dec_AND_node_2 S0 gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1012 D1 DEC_D1_NAND gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1013 D2 DEC_D2_NAND gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1014 DEC_D3_NAND S1 DEC_AND_NODE_4 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1015 vdd S0 DEC_D3_NAND vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1016 D2 DEC_D2_NAND vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1017 S0c S0 vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1018 DEC_D0_NAND S0c vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1019 D0 DEC_D0_NAND vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1020 D1 DEC_D1_NAND vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1021 DEC_AND_NODE_4 S0 gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1022 S1c S1 gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1023 DEC_D2_NAND S0c vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1024 D3 DEC_D3_NAND gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1025 vdd S1 DEC_D2_NAND vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1026 vdd S1c DEC_D0_NAND vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1027 DEC_D0_NAND S0c Dec_AND_node_1 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
C0 vdd D0 0.040884f
C1 DEC_D0_NAND Dec_AND_node_1 0.085282f
C2 S0 S1c 0.07308f
C3 vdd DEC_D0_NAND 0.094023f
C4 Dec_AND_node_1 S0c 0.088221f
C5 S1c gnd 0.055406f
C6 DEC_D2_NAND S0c 0.006448f
C7 vdd S0c 0.230788f
C8 D1 vdd 0.04098f
C9 Dec_AND_node_2 S1c 0.088221f
C10 S0 vdd 0.202099f
C11 S1 DEC_AND_NODE_4 0.088221f
C12 DEC_D3_NAND vdd 0.094059f
C13 Dec_AND_node_1 gnd 0.07683f
C14 DEC_D0_NAND D0 0.030251f
C15 DEC_D2_NAND gnd 0.157853f
C16 DEC_D2_NAND DEC_AND_NODE_3 0.085282f
C17 D1 DEC_D1_NAND 0.030251f
C18 vdd gnd 0.040225f
C19 vdd D3 0.04098f
C20 S1 S0c 0.511187f
C21 DEC_D2_NAND D2 0.030251f
C22 S0 DEC_D1_NAND 0.015311f
C23 vdd D2 0.04098f
C24 S0 S1 0.028532f
C25 DEC_D3_NAND S1 0.006448f
C26 DEC_D0_NAND S0c 0.006448f
C27 DEC_D1_NAND gnd 0.159401f
C28 S1 gnd 0.131827f
C29 S1 DEC_AND_NODE_3 0.089107f
C30 Dec_AND_node_2 DEC_D1_NAND 0.085282f
C31 S0 DEC_AND_NODE_4 0.089107f
C32 D0 gnd 0.051616f
C33 DEC_D3_NAND DEC_AND_NODE_4 0.085282f
C34 S1c Dec_AND_node_1 0.089107f
C35 DEC_D0_NAND gnd 0.145266f
C36 S0 S0c 0.043542f
C37 gnd DEC_AND_NODE_4 0.077062f
C38 vdd S1c 0.19269f
C39 gnd S0c 0.051616f
C40 D1 gnd 0.051616f
C41 S0 DEC_D3_NAND 0.015311f
C42 DEC_AND_NODE_3 S0c 0.088221f
C43 S0 gnd 0.092334f
C44 S1c DEC_D1_NAND 0.006448f
C45 DEC_D3_NAND gnd 0.157853f
C46 DEC_D3_NAND D3 0.030251f
C47 S1c S1 0.030251f
C48 vdd DEC_D2_NAND 0.094003f
C49 S0 Dec_AND_node_2 0.089107f
C50 gnd D3 0.051616f
C51 gnd DEC_AND_NODE_3 0.077196f
C52 S1c DEC_D0_NAND 0.015311f
C53 Dec_AND_node_2 gnd 0.077312f
C54 gnd D2 0.051616f
C55 DEC_D2_NAND S1 0.015311f
C56 vdd DEC_D1_NAND 0.094035f
C57 vdd S1 0.201098f
C58 S1c S0c 0.015985f
C59 DEC_AND_NODE_4 0 0.248064f **FLOATING
C60 D3 0 0.114466f **FLOATING
C61 DEC_D3_NAND 0 0.516966f **FLOATING
C62 DEC_AND_NODE_3 0 0.248064f **FLOATING
C63 D2 0 0.114466f **FLOATING
C64 DEC_D2_NAND 0 0.52029f **FLOATING
C65 Dec_AND_node_2 0 0.248064f **FLOATING
C66 S1 0 2.76414f **FLOATING
C67 D1 0 0.104663f **FLOATING
C68 DEC_D1_NAND 0 0.513722f **FLOATING
C69 S0 0 7.918251f **FLOATING
C70 gnd 0 8.80989f **FLOATING
C71 Dec_AND_node_1 0 0.248064f **FLOATING
C72 D0 0 0.075352f **FLOATING
C73 DEC_D0_NAND 0 0.511796f **FLOATING
C74 S1c 0 4.36861f **FLOATING
C75 S0c 0 5.09312f **FLOATING
C76 vdd 0 14.7771f **FLOATING
