magic
tech scmos
timestamp 1701340679
<< nwell >>
rect 157 388 218 405
rect 230 373 276 392
rect 156 270 217 287
rect 229 254 275 273
rect 2 234 86 253
rect 155 166 216 183
rect 230 150 276 169
rect 155 70 216 87
rect 228 54 275 73
<< ntransistor >>
rect 177 365 182 370
rect 200 365 205 370
rect 256 358 261 363
rect 176 247 181 252
rect 199 247 204 252
rect 28 219 33 224
rect 66 219 71 224
rect 255 239 260 244
rect 175 143 180 148
rect 198 143 203 148
rect 256 135 261 140
rect 175 47 180 52
rect 198 47 203 52
rect 255 39 260 44
<< ptransistor >>
rect 177 394 182 399
rect 200 394 205 399
rect 256 380 261 385
rect 176 276 181 281
rect 199 276 204 281
rect 255 261 260 266
rect 28 241 33 246
rect 66 241 71 246
rect 175 172 180 177
rect 198 172 203 177
rect 256 157 261 162
rect 175 76 180 81
rect 198 76 203 81
rect 255 61 260 66
<< ndiffusion >>
rect 175 365 177 370
rect 182 365 184 370
rect 198 365 200 370
rect 205 365 207 370
rect 254 358 256 363
rect 261 358 264 363
rect 174 247 176 252
rect 181 247 183 252
rect 197 247 199 252
rect 204 247 206 252
rect 26 219 28 224
rect 33 219 36 224
rect 64 219 66 224
rect 71 219 74 224
rect 253 239 255 244
rect 260 239 263 244
rect 173 143 175 148
rect 180 143 182 148
rect 196 143 198 148
rect 203 143 205 148
rect 254 135 256 140
rect 261 135 264 140
rect 173 47 175 52
rect 180 47 182 52
rect 196 47 198 52
rect 203 47 205 52
rect 253 39 255 44
rect 260 39 263 44
<< pdiffusion >>
rect 175 394 177 399
rect 182 394 189 399
rect 194 394 200 399
rect 205 394 207 399
rect 254 380 256 385
rect 261 380 264 385
rect 174 276 176 281
rect 181 276 188 281
rect 193 276 199 281
rect 204 276 206 281
rect 253 261 255 266
rect 260 261 263 266
rect 26 241 28 246
rect 33 241 36 246
rect 64 241 66 246
rect 71 241 74 246
rect 173 172 175 177
rect 180 172 187 177
rect 192 172 198 177
rect 203 172 205 177
rect 254 157 256 162
rect 261 157 264 162
rect 173 76 175 81
rect 180 76 187 81
rect 192 76 198 81
rect 203 76 205 81
rect 253 61 255 66
rect 260 61 263 66
<< ndcontact >>
rect 170 365 175 370
rect 184 365 188 370
rect 194 365 198 370
rect 207 365 212 370
rect 249 358 254 363
rect 264 358 269 363
rect 169 247 174 252
rect 183 247 187 252
rect 193 247 197 252
rect 206 247 211 252
rect 21 219 26 224
rect 36 219 41 224
rect 59 219 64 224
rect 74 219 79 224
rect 248 239 253 244
rect 263 239 268 244
rect 168 143 173 148
rect 182 143 186 148
rect 192 143 196 148
rect 205 143 210 148
rect 249 135 254 140
rect 264 135 269 140
rect 168 47 173 52
rect 182 47 186 52
rect 192 47 196 52
rect 205 47 210 52
rect 248 39 253 44
rect 263 39 268 44
<< pdcontact >>
rect 170 394 175 399
rect 189 394 194 399
rect 207 394 212 399
rect 249 380 254 385
rect 264 380 269 385
rect 169 276 174 281
rect 188 276 193 281
rect 206 276 211 281
rect 248 261 253 266
rect 263 261 268 266
rect 21 241 26 246
rect 36 241 41 246
rect 59 241 64 246
rect 74 241 79 246
rect 168 172 173 177
rect 187 172 192 177
rect 205 172 210 177
rect 249 157 254 162
rect 264 157 269 162
rect 168 76 173 81
rect 187 76 192 81
rect 205 76 210 81
rect 248 61 253 66
rect 263 61 268 66
<< nsubstratencontact >>
rect 161 394 166 399
rect 237 380 242 385
rect 160 276 165 281
rect 236 261 241 266
rect 9 241 14 246
rect 159 172 164 177
rect 237 157 242 162
rect 159 76 164 81
rect 236 61 241 66
<< polysilicon >>
rect 177 399 182 413
rect 200 399 205 413
rect 177 370 182 394
rect 200 370 205 394
rect 256 385 261 388
rect 256 371 261 380
rect 257 367 261 371
rect 177 346 182 365
rect 200 346 205 365
rect 256 363 261 367
rect 256 354 261 358
rect 176 281 181 295
rect 199 281 204 295
rect 176 252 181 276
rect 199 252 204 276
rect 255 266 260 269
rect 255 252 260 261
rect 28 246 33 249
rect 66 246 71 249
rect 256 248 260 252
rect 28 232 33 241
rect 66 232 71 241
rect 29 228 33 232
rect 67 228 71 232
rect 28 224 33 228
rect 66 224 71 228
rect 176 228 181 247
rect 199 228 204 247
rect 255 244 260 248
rect 255 234 260 239
rect 28 214 33 219
rect 66 214 71 219
rect 175 177 180 191
rect 198 177 203 191
rect 175 148 180 172
rect 198 148 203 172
rect 256 162 261 165
rect 256 148 261 157
rect 257 144 261 148
rect 175 124 180 143
rect 198 124 203 143
rect 256 140 261 144
rect 256 130 261 135
rect 175 81 180 95
rect 198 81 203 95
rect 175 52 180 76
rect 198 52 203 76
rect 255 66 260 69
rect 255 52 260 61
rect 256 48 260 52
rect 175 28 180 47
rect 198 28 203 47
rect 255 44 260 48
rect 255 34 260 39
<< polycontact >>
rect 252 367 257 371
rect 177 340 182 346
rect 200 340 205 346
rect 251 248 256 252
rect 24 228 29 232
rect 62 228 67 232
rect 176 222 181 228
rect 199 222 204 228
rect 252 144 257 148
rect 175 118 180 124
rect 198 118 203 124
rect 251 48 256 52
rect 175 22 180 28
rect 198 22 203 28
<< metal1 >>
rect 83 410 88 412
rect 209 410 312 411
rect 83 407 313 410
rect 83 406 212 407
rect 83 258 88 406
rect 161 405 212 406
rect 161 399 166 405
rect 170 399 175 405
rect 207 399 212 405
rect 232 397 236 407
rect 305 397 313 407
rect 189 384 194 394
rect 230 392 313 397
rect 184 380 194 384
rect 237 385 242 392
rect 249 385 254 392
rect 184 376 188 380
rect 184 373 225 376
rect 184 370 188 373
rect 222 370 225 373
rect 264 371 269 380
rect 229 370 252 371
rect 167 354 170 368
rect 212 365 214 368
rect 222 367 252 370
rect 264 367 272 371
rect 222 366 249 367
rect 194 362 197 365
rect 211 354 214 365
rect 264 363 269 367
rect 249 354 254 358
rect 167 349 214 354
rect 246 349 278 354
rect 2 253 88 258
rect 9 246 14 253
rect 21 246 26 253
rect 59 246 64 253
rect 22 228 24 232
rect 22 227 23 228
rect 36 224 41 241
rect 74 232 79 241
rect 59 228 62 232
rect 74 227 77 232
rect 74 224 79 227
rect 21 215 26 219
rect 59 217 64 219
rect 46 215 65 217
rect 10 214 91 215
rect 10 210 49 214
rect 62 212 91 214
rect 64 210 91 212
rect 10 5 16 210
rect 54 106 58 205
rect 100 118 108 326
rect 208 292 239 293
rect 160 289 239 292
rect 160 287 211 289
rect 160 281 165 287
rect 169 281 174 287
rect 206 281 211 287
rect 231 278 235 289
rect 305 278 313 392
rect 188 266 193 276
rect 229 273 313 278
rect 183 262 193 266
rect 236 266 241 273
rect 183 258 187 262
rect 248 266 253 273
rect 286 272 300 273
rect 183 255 224 258
rect 183 252 187 255
rect 221 252 224 255
rect 263 252 268 261
rect 166 236 169 250
rect 211 247 213 250
rect 221 248 251 252
rect 263 248 280 252
rect 193 244 196 247
rect 210 236 213 247
rect 263 244 268 248
rect 166 231 213 236
rect 248 235 253 239
rect 244 230 274 235
rect 176 219 181 222
rect 198 219 204 222
rect 207 188 238 189
rect 159 185 238 188
rect 159 183 210 185
rect 159 177 164 183
rect 168 177 173 183
rect 205 177 210 183
rect 230 174 234 185
rect 305 174 313 273
rect 187 162 192 172
rect 230 169 313 174
rect 182 158 192 162
rect 237 162 242 169
rect 182 154 186 158
rect 249 162 254 169
rect 182 151 223 154
rect 182 148 186 151
rect 220 148 223 151
rect 264 148 269 157
rect 165 132 168 146
rect 210 143 212 146
rect 220 144 252 148
rect 264 144 284 148
rect 192 140 195 143
rect 209 132 212 143
rect 264 140 269 144
rect 165 127 212 132
rect 249 131 254 135
rect 243 126 270 131
rect 100 113 180 118
rect 198 106 203 118
rect 54 100 203 106
rect 145 23 149 100
rect 207 92 238 93
rect 159 89 238 92
rect 159 87 210 89
rect 159 81 164 87
rect 168 81 173 87
rect 205 81 210 87
rect 230 78 234 89
rect 305 78 313 169
rect 187 66 192 76
rect 228 73 313 78
rect 182 62 192 66
rect 236 66 241 73
rect 182 58 186 62
rect 248 66 253 73
rect 182 55 223 58
rect 182 52 186 55
rect 220 52 223 55
rect 263 52 268 61
rect 165 36 168 50
rect 210 47 212 50
rect 220 48 251 52
rect 263 48 283 52
rect 192 44 195 47
rect 209 36 212 47
rect 263 44 268 48
rect 165 31 212 36
rect 248 35 253 39
rect 269 35 278 36
rect 244 30 278 35
rect 269 29 278 30
rect 145 22 175 23
rect 145 19 180 22
rect 271 5 277 29
rect 10 0 277 5
<< m2contact >>
rect 192 357 197 362
rect 239 348 246 354
rect 100 326 108 334
rect 177 333 182 340
rect 200 334 205 340
rect 17 227 22 232
rect 41 227 47 232
rect 54 227 59 232
rect 77 227 85 232
rect 53 205 59 210
rect 191 239 196 244
rect 236 230 244 235
rect 176 214 181 219
rect 198 213 204 219
rect 190 135 195 140
rect 235 126 243 132
rect 190 39 195 44
rect 236 29 244 35
rect 198 15 203 22
<< metal2 >>
rect 197 357 223 360
rect 218 353 223 357
rect 218 349 239 353
rect 218 348 230 349
rect 45 326 100 331
rect 177 331 182 333
rect 108 326 182 331
rect 45 234 50 326
rect 200 316 205 334
rect 132 309 205 316
rect 45 232 49 234
rect 132 232 139 309
rect 196 239 219 242
rect 0 227 17 232
rect 47 227 49 232
rect 85 227 139 232
rect 214 235 219 239
rect 223 235 228 348
rect 214 230 236 235
rect 0 201 6 227
rect 54 210 58 227
rect 132 215 139 227
rect 132 214 176 215
rect 132 208 181 214
rect 198 201 204 213
rect 0 197 204 201
rect 0 196 6 197
rect 40 15 44 197
rect 195 135 219 138
rect 214 131 219 135
rect 223 131 228 230
rect 214 126 235 131
rect 195 39 218 42
rect 214 35 218 39
rect 223 35 228 126
rect 214 30 236 35
rect 40 12 203 15
rect 198 11 203 12
<< labels >>
rlabel metal1 38 230 38 230 1 S0c
rlabel metal1 23 230 23 230 1 S0
rlabel metal1 61 231 61 231 1 S1
rlabel metal1 277 250 277 250 1 D1
rlabel metal1 271 369 271 369 1 D0
rlabel metal1 279 50 279 50 1 D3
rlabel metal1 188 33 188 33 1 DEC_AND_NODE_4
rlabel metal1 188 56 188 56 1 DEC_D3_NAND
rlabel metal1 280 146 280 146 1 D2
rlabel metal1 189 129 189 129 1 DEC_AND_NODE_3
rlabel metal1 189 152 189 152 1 DEC_D2_NAND
rlabel metal1 191 233 191 233 1 Dec_AND_node_2
rlabel metal1 192 256 192 256 1 DEC_D1_NAND
rlabel metal1 187 375 187 375 1 DEC_D0_NAND
rlabel metal1 192 352 192 352 1 Dec_AND_node_1
rlabel m2contact 80 230 80 230 1 S1c
rlabel metal1 80 212 80 212 1 gnd
rlabel metal1 56 256 56 256 1 vdd
<< end >>
