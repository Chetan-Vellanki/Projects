magic
tech scmos
timestamp 1701348530
<< nwell >>
rect 465 566 525 583
rect 539 550 585 569
rect 600 566 661 583
rect 675 550 721 569
rect 746 568 807 585
rect 821 552 867 571
rect 894 568 954 585
rect 968 552 1014 571
rect 1105 567 1166 584
rect 1180 551 1226 570
rect 1241 567 1302 584
rect 1316 551 1362 570
rect 1387 569 1448 586
rect 1462 553 1508 572
rect 1534 569 1595 586
rect 1609 553 1655 572
rect 464 458 525 475
rect 539 442 585 461
rect 608 458 669 475
rect 683 442 729 461
rect 757 460 818 477
rect 832 444 878 463
rect 902 461 963 478
rect 977 445 1023 464
rect 157 388 218 405
rect 230 373 276 392
rect 156 270 217 287
rect 229 254 275 273
rect 2 234 86 253
rect 155 166 216 183
rect 230 150 276 169
rect 155 70 216 87
rect 228 54 275 73
<< ntransistor >>
rect 484 543 489 548
rect 507 543 512 548
rect 620 543 625 548
rect 643 543 648 548
rect 766 545 771 550
rect 789 545 794 550
rect 565 535 570 540
rect 701 535 706 540
rect 913 545 918 550
rect 936 545 941 550
rect 847 537 852 542
rect 1125 544 1130 549
rect 1148 544 1153 549
rect 994 537 999 542
rect 1261 544 1266 549
rect 1284 544 1289 549
rect 1407 546 1412 551
rect 1430 546 1435 551
rect 1206 536 1211 541
rect 1342 536 1347 541
rect 1554 546 1559 551
rect 1577 546 1582 551
rect 1488 538 1493 543
rect 1635 538 1640 543
rect 484 435 489 440
rect 507 435 512 440
rect 628 435 633 440
rect 651 435 656 440
rect 777 437 782 442
rect 800 437 805 442
rect 922 438 927 443
rect 945 438 950 443
rect 565 427 570 432
rect 709 427 714 432
rect 858 429 863 434
rect 1003 430 1008 435
rect 177 365 182 370
rect 200 365 205 370
rect 256 358 261 363
rect 176 247 181 252
rect 199 247 204 252
rect 28 219 33 224
rect 66 219 71 224
rect 255 239 260 244
rect 175 143 180 148
rect 198 143 203 148
rect 256 135 261 140
rect 175 47 180 52
rect 198 47 203 52
rect 255 39 260 44
<< ptransistor >>
rect 484 572 489 577
rect 507 572 512 577
rect 620 572 625 577
rect 643 572 648 577
rect 766 574 771 579
rect 789 574 794 579
rect 913 574 918 579
rect 936 574 941 579
rect 565 557 570 562
rect 701 557 706 562
rect 847 559 852 564
rect 1125 573 1130 578
rect 1148 573 1153 578
rect 1261 573 1266 578
rect 1284 573 1289 578
rect 1407 575 1412 580
rect 1430 575 1435 580
rect 1554 575 1559 580
rect 1577 575 1582 580
rect 994 559 999 564
rect 1206 558 1211 563
rect 1342 558 1347 563
rect 1488 560 1493 565
rect 1635 560 1640 565
rect 484 464 489 469
rect 507 464 512 469
rect 628 464 633 469
rect 651 464 656 469
rect 777 466 782 471
rect 800 466 805 471
rect 922 467 927 472
rect 945 467 950 472
rect 565 449 570 454
rect 709 449 714 454
rect 858 451 863 456
rect 1003 452 1008 457
rect 177 394 182 399
rect 200 394 205 399
rect 256 380 261 385
rect 176 276 181 281
rect 199 276 204 281
rect 255 261 260 266
rect 28 241 33 246
rect 66 241 71 246
rect 175 172 180 177
rect 198 172 203 177
rect 256 157 261 162
rect 175 76 180 81
rect 198 76 203 81
rect 255 61 260 66
<< ndiffusion >>
rect 482 543 484 548
rect 489 543 491 548
rect 505 543 507 548
rect 512 543 514 548
rect 618 543 620 548
rect 625 543 627 548
rect 641 543 643 548
rect 648 543 650 548
rect 764 545 766 550
rect 771 545 773 550
rect 787 545 789 550
rect 794 545 796 550
rect 563 535 565 540
rect 570 535 573 540
rect 699 535 701 540
rect 706 535 709 540
rect 911 545 913 550
rect 918 545 920 550
rect 934 545 936 550
rect 941 545 943 550
rect 845 537 847 542
rect 852 537 855 542
rect 1123 544 1125 549
rect 1130 544 1132 549
rect 1146 544 1148 549
rect 1153 544 1155 549
rect 992 537 994 542
rect 999 537 1002 542
rect 1259 544 1261 549
rect 1266 544 1268 549
rect 1282 544 1284 549
rect 1289 544 1291 549
rect 1405 546 1407 551
rect 1412 546 1414 551
rect 1428 546 1430 551
rect 1435 546 1437 551
rect 1204 536 1206 541
rect 1211 536 1214 541
rect 1340 536 1342 541
rect 1347 536 1350 541
rect 1552 546 1554 551
rect 1559 546 1561 551
rect 1575 546 1577 551
rect 1582 546 1584 551
rect 1486 538 1488 543
rect 1493 538 1496 543
rect 1633 538 1635 543
rect 1640 538 1643 543
rect 482 435 484 440
rect 489 435 491 440
rect 505 435 507 440
rect 512 435 514 440
rect 626 435 628 440
rect 633 435 635 440
rect 649 435 651 440
rect 656 435 658 440
rect 775 437 777 442
rect 782 437 784 442
rect 798 437 800 442
rect 805 437 807 442
rect 920 438 922 443
rect 927 438 929 443
rect 943 438 945 443
rect 950 438 952 443
rect 563 427 565 432
rect 570 427 573 432
rect 707 427 709 432
rect 714 427 717 432
rect 856 429 858 434
rect 863 429 866 434
rect 1001 430 1003 435
rect 1008 430 1011 435
rect 175 365 177 370
rect 182 365 184 370
rect 198 365 200 370
rect 205 365 207 370
rect 254 358 256 363
rect 261 358 264 363
rect 174 247 176 252
rect 181 247 183 252
rect 197 247 199 252
rect 204 247 206 252
rect 26 219 28 224
rect 33 219 36 224
rect 64 219 66 224
rect 71 219 74 224
rect 253 239 255 244
rect 260 239 263 244
rect 173 143 175 148
rect 180 143 182 148
rect 196 143 198 148
rect 203 143 205 148
rect 254 135 256 140
rect 261 135 264 140
rect 173 47 175 52
rect 180 47 182 52
rect 196 47 198 52
rect 203 47 205 52
rect 253 39 255 44
rect 260 39 263 44
<< pdiffusion >>
rect 482 572 484 577
rect 489 572 496 577
rect 501 572 507 577
rect 512 572 514 577
rect 618 572 620 577
rect 625 572 632 577
rect 637 572 643 577
rect 648 572 650 577
rect 764 574 766 579
rect 771 574 778 579
rect 783 574 789 579
rect 794 574 796 579
rect 911 574 913 579
rect 918 574 925 579
rect 930 574 936 579
rect 941 574 943 579
rect 563 557 565 562
rect 570 557 573 562
rect 699 557 701 562
rect 706 557 709 562
rect 845 559 847 564
rect 852 559 855 564
rect 1123 573 1125 578
rect 1130 573 1137 578
rect 1142 573 1148 578
rect 1153 573 1155 578
rect 1259 573 1261 578
rect 1266 573 1273 578
rect 1278 573 1284 578
rect 1289 573 1291 578
rect 1405 575 1407 580
rect 1412 575 1419 580
rect 1424 575 1430 580
rect 1435 575 1437 580
rect 1552 575 1554 580
rect 1559 575 1566 580
rect 1571 575 1577 580
rect 1582 575 1584 580
rect 992 559 994 564
rect 999 559 1002 564
rect 1204 558 1206 563
rect 1211 558 1214 563
rect 1340 558 1342 563
rect 1347 558 1350 563
rect 1486 560 1488 565
rect 1493 560 1496 565
rect 1633 560 1635 565
rect 1640 560 1643 565
rect 482 464 484 469
rect 489 464 496 469
rect 501 464 507 469
rect 512 464 514 469
rect 626 464 628 469
rect 633 464 640 469
rect 645 464 651 469
rect 656 464 658 469
rect 775 466 777 471
rect 782 466 789 471
rect 794 466 800 471
rect 805 466 807 471
rect 920 467 922 472
rect 927 467 934 472
rect 939 467 945 472
rect 950 467 952 472
rect 563 449 565 454
rect 570 449 573 454
rect 707 449 709 454
rect 714 449 717 454
rect 856 451 858 456
rect 863 451 866 456
rect 1001 452 1003 457
rect 1008 452 1011 457
rect 175 394 177 399
rect 182 394 189 399
rect 194 394 200 399
rect 205 394 207 399
rect 254 380 256 385
rect 261 380 264 385
rect 174 276 176 281
rect 181 276 188 281
rect 193 276 199 281
rect 204 276 206 281
rect 253 261 255 266
rect 260 261 263 266
rect 26 241 28 246
rect 33 241 36 246
rect 64 241 66 246
rect 71 241 74 246
rect 173 172 175 177
rect 180 172 187 177
rect 192 172 198 177
rect 203 172 205 177
rect 254 157 256 162
rect 261 157 264 162
rect 173 76 175 81
rect 180 76 187 81
rect 192 76 198 81
rect 203 76 205 81
rect 253 61 255 66
rect 260 61 263 66
<< ndcontact >>
rect 477 543 482 548
rect 491 543 495 548
rect 501 543 505 548
rect 514 543 519 548
rect 613 543 618 548
rect 627 543 631 548
rect 637 543 641 548
rect 650 543 655 548
rect 759 545 764 550
rect 773 545 777 550
rect 783 545 787 550
rect 796 545 801 550
rect 558 535 563 540
rect 573 535 578 540
rect 694 535 699 540
rect 709 535 714 540
rect 906 545 911 550
rect 920 545 924 550
rect 930 545 934 550
rect 943 545 948 550
rect 840 537 845 542
rect 855 537 860 542
rect 1118 544 1123 549
rect 1132 544 1136 549
rect 1142 544 1146 549
rect 1155 544 1160 549
rect 987 537 992 542
rect 1002 537 1007 542
rect 1254 544 1259 549
rect 1268 544 1272 549
rect 1278 544 1282 549
rect 1291 544 1296 549
rect 1400 546 1405 551
rect 1414 546 1418 551
rect 1424 546 1428 551
rect 1437 546 1442 551
rect 1199 536 1204 541
rect 1214 536 1219 541
rect 1335 536 1340 541
rect 1350 536 1355 541
rect 1547 546 1552 551
rect 1561 546 1565 551
rect 1571 546 1575 551
rect 1584 546 1589 551
rect 1481 538 1486 543
rect 1496 538 1501 543
rect 1628 538 1633 543
rect 1643 538 1648 543
rect 477 435 482 440
rect 491 435 495 440
rect 501 435 505 440
rect 514 435 519 440
rect 621 435 626 440
rect 635 435 639 440
rect 645 435 649 440
rect 658 435 663 440
rect 770 437 775 442
rect 784 437 788 442
rect 794 437 798 442
rect 807 437 812 442
rect 915 438 920 443
rect 929 438 933 443
rect 939 438 943 443
rect 952 438 957 443
rect 558 427 563 432
rect 573 427 578 432
rect 702 427 707 432
rect 717 427 722 432
rect 851 429 856 434
rect 866 429 871 434
rect 996 430 1001 435
rect 1011 430 1016 435
rect 170 365 175 370
rect 184 365 188 370
rect 194 365 198 370
rect 207 365 212 370
rect 249 358 254 363
rect 264 358 269 363
rect 169 247 174 252
rect 183 247 187 252
rect 193 247 197 252
rect 206 247 211 252
rect 21 219 26 224
rect 36 219 41 224
rect 59 219 64 224
rect 74 219 79 224
rect 248 239 253 244
rect 263 239 268 244
rect 168 143 173 148
rect 182 143 186 148
rect 192 143 196 148
rect 205 143 210 148
rect 249 135 254 140
rect 264 135 269 140
rect 168 47 173 52
rect 182 47 186 52
rect 192 47 196 52
rect 205 47 210 52
rect 248 39 253 44
rect 263 39 268 44
<< pdcontact >>
rect 477 572 482 577
rect 496 572 501 577
rect 514 572 519 577
rect 613 572 618 577
rect 632 572 637 577
rect 650 572 655 577
rect 759 574 764 579
rect 778 574 783 579
rect 796 574 801 579
rect 906 574 911 579
rect 925 574 930 579
rect 943 574 948 579
rect 558 557 563 562
rect 573 557 578 562
rect 694 557 699 562
rect 709 557 714 562
rect 840 559 845 564
rect 855 559 860 564
rect 1118 573 1123 578
rect 1137 573 1142 578
rect 1155 573 1160 578
rect 1254 573 1259 578
rect 1273 573 1278 578
rect 1291 573 1296 578
rect 1400 575 1405 580
rect 1419 575 1424 580
rect 1437 575 1442 580
rect 1547 575 1552 580
rect 1566 575 1571 580
rect 1584 575 1589 580
rect 987 559 992 564
rect 1002 559 1007 564
rect 1199 558 1204 563
rect 1214 558 1219 563
rect 1335 558 1340 563
rect 1350 558 1355 563
rect 1481 560 1486 565
rect 1496 560 1501 565
rect 1628 560 1633 565
rect 1643 560 1648 565
rect 477 464 482 469
rect 496 464 501 469
rect 514 464 519 469
rect 621 464 626 469
rect 640 464 645 469
rect 658 464 663 469
rect 770 466 775 471
rect 789 466 794 471
rect 807 466 812 471
rect 915 467 920 472
rect 934 467 939 472
rect 952 467 957 472
rect 558 449 563 454
rect 573 449 578 454
rect 702 449 707 454
rect 717 449 722 454
rect 851 451 856 456
rect 866 451 871 456
rect 996 452 1001 457
rect 1011 452 1016 457
rect 170 394 175 399
rect 189 394 194 399
rect 207 394 212 399
rect 249 380 254 385
rect 264 380 269 385
rect 169 276 174 281
rect 188 276 193 281
rect 206 276 211 281
rect 248 261 253 266
rect 263 261 268 266
rect 21 241 26 246
rect 36 241 41 246
rect 59 241 64 246
rect 74 241 79 246
rect 168 172 173 177
rect 187 172 192 177
rect 205 172 210 177
rect 249 157 254 162
rect 264 157 269 162
rect 168 76 173 81
rect 187 76 192 81
rect 205 76 210 81
rect 248 61 253 66
rect 263 61 268 66
<< nsubstratencontact >>
rect 468 572 473 577
rect 604 572 609 577
rect 751 574 755 579
rect 897 574 902 579
rect 546 557 551 562
rect 682 557 687 562
rect 828 559 833 564
rect 1109 573 1114 578
rect 1245 573 1250 578
rect 1391 575 1396 580
rect 1538 575 1543 580
rect 975 559 980 564
rect 1187 558 1192 563
rect 1323 558 1328 563
rect 1469 560 1474 565
rect 1616 560 1621 565
rect 468 464 473 469
rect 612 464 617 469
rect 761 466 766 471
rect 906 467 911 472
rect 546 449 551 454
rect 690 449 695 454
rect 839 451 844 456
rect 984 452 989 457
rect 161 394 166 399
rect 237 380 242 385
rect 160 276 165 281
rect 236 261 241 266
rect 9 241 14 246
rect 159 172 164 177
rect 237 157 242 162
rect 159 76 164 81
rect 236 61 241 66
<< polysilicon >>
rect 484 577 489 591
rect 507 577 512 591
rect 620 577 625 591
rect 643 577 648 591
rect 766 579 771 593
rect 789 579 794 593
rect 913 579 918 593
rect 936 579 941 593
rect 1125 578 1130 592
rect 1148 578 1153 592
rect 1261 578 1266 592
rect 1284 578 1289 592
rect 1407 580 1412 594
rect 1430 580 1435 594
rect 1554 580 1559 594
rect 1577 580 1582 594
rect 484 548 489 572
rect 507 548 512 572
rect 565 562 570 565
rect 565 548 570 557
rect 620 548 625 572
rect 643 548 648 572
rect 701 562 706 565
rect 701 548 706 557
rect 766 550 771 574
rect 789 550 794 574
rect 847 564 852 567
rect 847 550 852 559
rect 913 550 918 574
rect 936 550 941 574
rect 994 564 999 567
rect 994 550 999 559
rect 566 544 570 548
rect 484 524 489 543
rect 507 524 512 543
rect 565 540 570 544
rect 702 544 706 548
rect 848 546 852 550
rect 565 530 570 535
rect 620 524 625 543
rect 643 524 648 543
rect 701 540 706 544
rect 701 530 706 535
rect 766 526 771 545
rect 789 526 794 545
rect 847 542 852 546
rect 995 546 999 550
rect 1125 549 1130 573
rect 1148 549 1153 573
rect 1206 563 1211 566
rect 1206 549 1211 558
rect 1261 549 1266 573
rect 1284 549 1289 573
rect 1342 563 1347 566
rect 1342 549 1347 558
rect 1407 551 1412 575
rect 1430 551 1435 575
rect 1488 565 1493 568
rect 1488 551 1493 560
rect 1554 551 1559 575
rect 1577 551 1582 575
rect 1635 565 1640 568
rect 1635 551 1640 560
rect 847 532 852 537
rect 913 526 918 545
rect 936 526 941 545
rect 994 542 999 546
rect 1207 545 1211 549
rect 994 532 999 537
rect 1125 525 1130 544
rect 1148 525 1153 544
rect 1206 541 1211 545
rect 1343 545 1347 549
rect 1489 547 1493 551
rect 1206 531 1211 536
rect 1261 525 1266 544
rect 1284 525 1289 544
rect 1342 541 1347 545
rect 1342 531 1347 536
rect 1407 527 1412 546
rect 1430 527 1435 546
rect 1488 543 1493 547
rect 1636 547 1640 551
rect 1488 533 1493 538
rect 1554 527 1559 546
rect 1577 527 1582 546
rect 1635 543 1640 547
rect 1635 533 1640 538
rect 484 469 489 483
rect 507 469 512 483
rect 628 469 633 483
rect 651 469 656 483
rect 777 471 782 485
rect 800 471 805 485
rect 922 472 927 486
rect 945 472 950 486
rect 484 440 489 464
rect 507 440 512 464
rect 565 454 570 457
rect 565 440 570 449
rect 628 440 633 464
rect 651 440 656 464
rect 709 454 714 457
rect 709 440 714 449
rect 777 442 782 466
rect 800 442 805 466
rect 858 456 863 459
rect 858 442 863 451
rect 922 443 927 467
rect 945 443 950 467
rect 1003 457 1008 460
rect 1003 443 1008 452
rect 566 436 570 440
rect 484 416 489 435
rect 177 399 182 413
rect 200 399 205 413
rect 507 416 512 435
rect 565 432 570 436
rect 710 436 714 440
rect 859 438 863 442
rect 1004 439 1008 443
rect 565 422 570 427
rect 628 416 633 435
rect 651 416 656 435
rect 709 432 714 436
rect 709 422 714 427
rect 777 418 782 437
rect 800 418 805 437
rect 858 434 863 438
rect 858 424 863 429
rect 922 419 927 438
rect 945 419 950 438
rect 1003 435 1008 439
rect 1003 425 1008 430
rect 177 370 182 394
rect 200 370 205 394
rect 256 385 261 388
rect 256 371 261 380
rect 257 367 261 371
rect 177 346 182 365
rect 200 346 205 365
rect 256 363 261 367
rect 256 354 261 358
rect 176 281 181 295
rect 199 281 204 295
rect 176 252 181 276
rect 199 252 204 276
rect 255 266 260 269
rect 255 252 260 261
rect 28 246 33 249
rect 66 246 71 249
rect 256 248 260 252
rect 28 232 33 241
rect 66 232 71 241
rect 29 228 33 232
rect 67 228 71 232
rect 28 224 33 228
rect 66 224 71 228
rect 176 228 181 247
rect 199 228 204 247
rect 255 244 260 248
rect 255 234 260 239
rect 28 214 33 219
rect 66 214 71 219
rect 175 177 180 191
rect 198 177 203 191
rect 175 148 180 172
rect 198 148 203 172
rect 256 162 261 165
rect 256 148 261 157
rect 257 144 261 148
rect 175 124 180 143
rect 198 124 203 143
rect 256 140 261 144
rect 256 130 261 135
rect 175 81 180 95
rect 198 81 203 95
rect 175 52 180 76
rect 198 52 203 76
rect 255 66 260 69
rect 255 52 260 61
rect 256 48 260 52
rect 175 28 180 47
rect 198 28 203 47
rect 255 44 260 48
rect 255 34 260 39
<< polycontact >>
rect 561 544 566 548
rect 484 518 489 524
rect 697 544 702 548
rect 843 546 848 550
rect 507 518 512 524
rect 620 518 625 524
rect 643 518 648 524
rect 766 520 771 526
rect 990 546 995 550
rect 789 520 794 526
rect 913 520 918 526
rect 1202 545 1207 549
rect 936 520 941 526
rect 1125 519 1130 525
rect 1338 545 1343 549
rect 1484 547 1489 551
rect 1148 519 1153 525
rect 1261 519 1266 525
rect 1284 519 1289 525
rect 1407 521 1412 527
rect 1631 547 1636 551
rect 1430 521 1435 527
rect 1554 521 1559 527
rect 1577 521 1582 527
rect 561 436 566 440
rect 484 410 489 416
rect 705 436 710 440
rect 854 438 859 442
rect 999 439 1004 443
rect 507 410 512 416
rect 628 410 633 416
rect 651 410 656 416
rect 777 412 782 418
rect 800 412 805 418
rect 922 413 927 419
rect 945 413 950 419
rect 252 367 257 371
rect 177 340 182 346
rect 200 340 205 346
rect 251 248 256 252
rect 24 228 29 232
rect 62 228 67 232
rect 176 222 181 228
rect 199 222 204 228
rect 252 144 257 148
rect 175 118 180 124
rect 198 118 203 124
rect 251 48 256 52
rect 175 22 180 28
rect 198 22 203 28
<< metal1 >>
rect 730 641 1230 646
rect 730 621 736 641
rect 883 618 1378 624
rect 305 588 312 593
rect 1439 591 1539 592
rect 1586 591 1617 592
rect 798 590 898 591
rect 945 590 976 591
rect 1391 590 1617 591
rect 744 589 976 590
rect 1157 589 1188 590
rect 1293 589 1617 590
rect 516 588 547 589
rect 652 588 976 589
rect 1102 588 1617 589
rect 305 587 1442 588
rect 305 585 801 587
rect 305 583 519 585
rect 83 410 88 412
rect 305 411 312 583
rect 447 582 474 583
rect 447 482 455 582
rect 468 577 473 582
rect 477 577 482 583
rect 514 577 519 583
rect 539 584 655 585
rect 539 574 543 584
rect 604 583 655 584
rect 604 577 609 583
rect 496 562 501 572
rect 539 569 587 574
rect 613 577 618 583
rect 650 577 655 583
rect 675 574 679 585
rect 751 579 755 585
rect 759 579 764 585
rect 796 579 801 585
rect 821 576 825 587
rect 897 585 948 587
rect 897 579 902 585
rect 491 558 501 562
rect 546 562 551 569
rect 491 554 495 558
rect 558 562 563 569
rect 632 562 637 572
rect 675 569 723 574
rect 491 551 532 554
rect 491 548 495 551
rect 529 548 532 551
rect 573 548 578 557
rect 627 558 637 562
rect 682 562 687 569
rect 627 554 631 558
rect 694 562 699 569
rect 778 564 783 574
rect 821 571 869 576
rect 906 579 911 585
rect 943 579 948 585
rect 968 586 1442 587
rect 968 584 1160 586
rect 968 576 972 584
rect 1102 583 1115 584
rect 1109 578 1114 583
rect 627 551 668 554
rect 474 532 477 546
rect 519 543 521 546
rect 529 544 561 548
rect 573 544 592 548
rect 501 540 504 543
rect 518 532 521 543
rect 573 540 578 544
rect 627 548 631 551
rect 665 548 668 551
rect 709 548 714 557
rect 773 560 783 564
rect 828 564 833 571
rect 773 556 777 560
rect 840 564 845 571
rect 925 564 930 574
rect 968 571 1016 576
rect 1118 578 1123 584
rect 1155 578 1160 584
rect 1180 585 1296 586
rect 1180 575 1184 585
rect 1245 584 1296 585
rect 1245 578 1250 584
rect 773 553 814 556
rect 773 550 777 553
rect 811 550 814 553
rect 855 550 860 559
rect 920 560 930 564
rect 975 564 980 571
rect 920 556 924 560
rect 987 564 992 571
rect 1137 563 1142 573
rect 1180 570 1228 575
rect 1254 578 1259 584
rect 1291 578 1296 584
rect 1316 575 1320 586
rect 1391 580 1396 586
rect 1400 580 1405 586
rect 1437 580 1442 586
rect 1462 577 1466 588
rect 1538 586 1589 588
rect 1538 580 1543 586
rect 920 553 961 556
rect 474 527 521 532
rect 558 531 563 535
rect 610 532 613 546
rect 655 543 657 546
rect 665 544 697 548
rect 709 544 730 548
rect 637 540 640 543
rect 654 532 657 543
rect 709 540 714 544
rect 553 526 588 531
rect 610 527 657 532
rect 484 517 489 518
rect 507 517 512 518
rect 584 505 588 526
rect 694 531 699 535
rect 756 534 759 548
rect 801 545 803 548
rect 811 546 843 550
rect 855 546 876 550
rect 783 542 786 545
rect 800 534 803 545
rect 855 542 860 546
rect 920 550 924 553
rect 958 550 961 553
rect 1002 550 1007 559
rect 1132 559 1142 563
rect 1187 563 1192 570
rect 1132 555 1136 559
rect 1199 563 1204 570
rect 1273 563 1278 573
rect 1316 570 1364 575
rect 1132 552 1173 555
rect 689 530 724 531
rect 689 526 737 530
rect 756 529 803 534
rect 840 533 845 537
rect 903 534 906 548
rect 948 545 950 548
rect 958 546 990 550
rect 1002 546 1032 550
rect 930 542 933 545
rect 947 534 950 545
rect 1002 542 1007 546
rect 1132 549 1136 552
rect 1170 549 1173 552
rect 1214 549 1219 558
rect 1268 559 1278 563
rect 1323 563 1328 570
rect 1268 555 1272 559
rect 1335 563 1340 570
rect 1419 565 1424 575
rect 1462 572 1510 577
rect 1547 580 1552 586
rect 1584 580 1589 586
rect 1609 577 1613 588
rect 1268 552 1309 555
rect 1268 549 1272 552
rect 1306 549 1309 552
rect 1350 549 1355 558
rect 1414 561 1424 565
rect 1469 565 1474 572
rect 1414 557 1418 561
rect 1481 565 1486 572
rect 1566 565 1571 575
rect 1609 572 1657 577
rect 1414 554 1455 557
rect 1414 551 1418 554
rect 1452 551 1455 554
rect 1496 551 1501 560
rect 1561 561 1571 565
rect 1616 565 1621 572
rect 1561 557 1565 561
rect 1628 565 1633 572
rect 1561 554 1602 557
rect 1561 551 1565 554
rect 1599 551 1602 554
rect 1643 551 1648 560
rect 835 528 873 533
rect 903 529 950 534
rect 718 525 737 526
rect 620 517 625 518
rect 643 517 648 518
rect 728 505 735 525
rect 766 519 771 520
rect 789 519 794 520
rect 864 505 873 528
rect 987 533 992 537
rect 1115 533 1118 547
rect 1160 544 1162 547
rect 1170 545 1202 549
rect 1214 545 1222 549
rect 1142 541 1145 544
rect 1159 533 1162 544
rect 1214 541 1219 545
rect 982 528 1018 533
rect 1115 528 1162 533
rect 913 519 918 520
rect 936 519 941 520
rect 1009 505 1018 528
rect 1199 532 1204 536
rect 1251 533 1254 547
rect 1296 544 1298 547
rect 1306 545 1338 549
rect 1350 545 1358 549
rect 1278 541 1281 544
rect 1295 533 1298 544
rect 1350 541 1355 545
rect 1194 527 1229 532
rect 1251 528 1298 533
rect 1125 518 1130 519
rect 1148 518 1153 519
rect 1225 506 1229 527
rect 1335 532 1340 536
rect 1397 535 1400 549
rect 1442 546 1444 549
rect 1452 547 1484 551
rect 1496 547 1504 551
rect 1424 543 1427 546
rect 1441 535 1444 546
rect 1496 543 1501 547
rect 1330 531 1365 532
rect 1330 527 1378 531
rect 1397 530 1444 535
rect 1481 534 1486 538
rect 1544 535 1547 549
rect 1589 546 1591 549
rect 1599 547 1631 551
rect 1643 547 1651 551
rect 1571 543 1574 546
rect 1588 535 1591 546
rect 1643 543 1648 547
rect 1476 529 1514 534
rect 1544 530 1591 535
rect 1359 526 1378 527
rect 1261 518 1266 519
rect 1284 518 1289 519
rect 1369 506 1376 526
rect 1407 520 1412 521
rect 1430 520 1435 521
rect 1505 506 1514 529
rect 1628 534 1633 538
rect 1623 529 1659 534
rect 1554 520 1559 521
rect 1577 520 1582 521
rect 1650 506 1659 529
rect 1037 505 1045 506
rect 584 499 1045 505
rect 1225 501 1660 506
rect 1225 500 1635 501
rect 1037 488 1045 499
rect 1246 488 1255 500
rect 954 483 985 484
rect 809 482 985 483
rect 447 480 477 482
rect 685 481 985 482
rect 516 480 547 481
rect 660 480 985 481
rect 1036 480 1255 488
rect 447 479 957 480
rect 447 477 812 479
rect 821 478 957 479
rect 447 475 519 477
rect 538 475 663 477
rect 468 469 473 475
rect 477 469 482 475
rect 514 469 519 475
rect 539 466 543 475
rect 612 469 617 475
rect 496 454 501 464
rect 539 461 587 466
rect 621 469 626 475
rect 658 469 663 475
rect 683 466 687 477
rect 761 471 766 477
rect 770 471 775 477
rect 807 471 812 477
rect 832 468 836 478
rect 906 472 911 478
rect 491 450 501 454
rect 546 454 551 461
rect 491 446 495 450
rect 558 454 563 461
rect 640 454 645 464
rect 683 461 731 466
rect 491 443 532 446
rect 491 440 495 443
rect 529 440 532 443
rect 573 440 578 449
rect 635 450 645 454
rect 690 454 695 461
rect 635 446 639 450
rect 702 454 707 461
rect 789 456 794 466
rect 832 463 880 468
rect 915 472 920 478
rect 952 472 957 478
rect 977 469 981 480
rect 635 443 676 446
rect 474 424 477 438
rect 519 435 521 438
rect 529 436 561 440
rect 573 436 605 440
rect 501 432 504 435
rect 518 424 521 435
rect 573 432 578 436
rect 635 440 639 443
rect 673 440 676 443
rect 717 440 722 449
rect 784 452 794 456
rect 839 456 844 463
rect 784 448 788 452
rect 851 456 856 463
rect 934 457 939 467
rect 977 464 1025 469
rect 784 445 825 448
rect 784 442 788 445
rect 822 442 825 445
rect 866 442 871 451
rect 929 453 939 457
rect 984 457 989 464
rect 929 449 933 453
rect 996 457 1001 464
rect 929 446 970 449
rect 929 443 933 446
rect 967 443 970 446
rect 1011 443 1016 452
rect 474 419 521 424
rect 558 423 563 427
rect 618 424 621 438
rect 663 435 665 438
rect 673 436 705 440
rect 717 436 745 440
rect 645 432 648 435
rect 662 424 665 435
rect 717 432 722 436
rect 553 418 588 423
rect 618 419 665 424
rect 209 410 312 411
rect 83 407 313 410
rect 83 406 212 407
rect 83 258 88 406
rect 161 405 212 406
rect 161 399 166 405
rect 170 399 175 405
rect 207 399 212 405
rect 232 397 236 407
rect 305 397 313 407
rect 484 409 489 410
rect 507 409 512 410
rect 189 384 194 394
rect 230 392 313 397
rect 184 380 194 384
rect 237 385 242 392
rect 249 385 254 392
rect 184 376 188 380
rect 184 373 225 376
rect 184 370 188 373
rect 222 370 225 373
rect 264 371 269 380
rect 305 372 313 392
rect 580 394 589 418
rect 702 423 707 427
rect 767 426 770 440
rect 812 437 814 440
rect 822 438 854 442
rect 866 438 894 442
rect 794 434 797 437
rect 811 426 814 437
rect 866 434 871 438
rect 697 418 738 423
rect 767 421 814 426
rect 851 425 856 429
rect 912 427 915 441
rect 957 438 959 441
rect 967 439 999 443
rect 1011 439 1019 443
rect 939 435 942 438
rect 956 427 959 438
rect 1011 435 1016 439
rect 846 420 881 425
rect 912 422 959 427
rect 996 426 1001 430
rect 1020 426 1027 427
rect 991 421 1027 426
rect 628 409 633 410
rect 651 409 656 410
rect 730 394 737 418
rect 777 411 782 412
rect 800 411 805 412
rect 874 394 881 420
rect 922 411 927 413
rect 945 412 950 413
rect 1020 394 1027 421
rect 580 393 1027 394
rect 1037 393 1045 480
rect 1246 479 1255 480
rect 580 388 1045 393
rect 229 370 252 371
rect 167 354 170 368
rect 212 365 214 368
rect 222 367 252 370
rect 264 367 272 371
rect 222 366 249 367
rect 194 362 197 365
rect 211 354 214 365
rect 264 363 269 367
rect 306 367 312 372
rect 249 354 254 358
rect 167 349 214 354
rect 246 349 268 354
rect 261 348 268 349
rect 2 253 88 258
rect 305 353 313 367
rect 304 348 314 353
rect 9 246 14 253
rect 21 246 26 253
rect 59 246 64 253
rect 22 228 24 232
rect 22 227 23 228
rect 36 224 41 241
rect 74 232 79 241
rect 59 228 62 232
rect 74 227 77 232
rect 74 224 79 227
rect 21 215 26 219
rect 59 217 64 219
rect 46 215 65 217
rect 10 214 91 215
rect 10 210 49 214
rect 62 212 91 214
rect 64 210 91 212
rect 10 5 16 210
rect 54 106 58 205
rect 100 118 108 326
rect 208 292 239 293
rect 160 289 239 292
rect 160 287 211 289
rect 160 281 165 287
rect 169 281 174 287
rect 206 281 211 287
rect 231 278 235 289
rect 305 278 313 348
rect 547 353 556 355
rect 341 348 556 353
rect 547 319 556 348
rect 688 319 695 388
rect 730 386 737 388
rect 1020 387 1027 388
rect 547 313 696 319
rect 688 311 695 313
rect 188 266 193 276
rect 229 273 313 278
rect 183 262 193 266
rect 236 266 241 273
rect 183 258 187 262
rect 248 266 253 273
rect 286 272 300 273
rect 183 255 224 258
rect 183 252 187 255
rect 221 252 224 255
rect 263 252 268 261
rect 166 236 169 250
rect 211 247 213 250
rect 221 248 251 252
rect 263 248 280 252
rect 193 244 196 247
rect 210 236 213 247
rect 263 244 268 248
rect 166 231 213 236
rect 248 235 253 239
rect 244 230 274 235
rect 176 219 181 222
rect 198 219 204 222
rect 207 188 238 189
rect 159 185 238 188
rect 159 183 210 185
rect 159 177 164 183
rect 168 177 173 183
rect 205 177 210 183
rect 230 174 234 185
rect 305 174 313 273
rect 187 162 192 172
rect 230 169 313 174
rect 182 158 192 162
rect 237 162 242 169
rect 182 154 186 158
rect 249 162 254 169
rect 182 151 223 154
rect 182 148 186 151
rect 220 148 223 151
rect 264 148 269 157
rect 165 132 168 146
rect 210 143 212 146
rect 220 144 252 148
rect 264 144 284 148
rect 192 140 195 143
rect 209 132 212 143
rect 264 140 269 144
rect 165 127 212 132
rect 249 131 254 135
rect 243 126 270 131
rect 100 113 180 118
rect 198 106 203 118
rect 54 100 203 106
rect 145 23 149 100
rect 207 92 238 93
rect 159 89 238 92
rect 159 87 210 89
rect 159 81 164 87
rect 168 81 173 87
rect 205 81 210 87
rect 230 78 234 89
rect 305 78 313 169
rect 187 66 192 76
rect 228 73 313 78
rect 182 62 192 66
rect 236 66 241 73
rect 182 58 186 62
rect 248 66 253 73
rect 182 55 223 58
rect 182 52 186 55
rect 220 52 223 55
rect 263 52 268 61
rect 165 36 168 50
rect 210 47 212 50
rect 220 48 251 52
rect 263 48 417 52
rect 192 44 195 47
rect 209 36 212 47
rect 263 44 268 48
rect 165 31 212 36
rect 248 35 253 39
rect 269 35 277 36
rect 244 30 277 35
rect 269 29 277 30
rect 145 22 175 23
rect 145 19 180 22
rect 271 5 277 29
rect 10 0 277 5
<< m2contact >>
rect 1230 638 1240 647
rect 726 614 736 621
rect 874 618 883 624
rect 1378 615 1388 625
rect 499 535 504 540
rect 592 542 598 549
rect 546 525 553 532
rect 635 535 640 540
rect 730 543 736 550
rect 484 510 489 517
rect 507 510 512 517
rect 682 525 689 532
rect 781 537 786 542
rect 876 544 882 551
rect 828 527 835 534
rect 928 537 933 542
rect 1032 544 1039 552
rect 620 510 625 517
rect 643 510 648 517
rect 766 512 771 519
rect 789 512 794 519
rect 975 527 982 534
rect 1140 536 1145 541
rect 913 512 918 519
rect 936 512 941 519
rect 1187 526 1194 533
rect 1276 536 1281 541
rect 1125 511 1130 518
rect 1148 511 1153 518
rect 1323 526 1330 533
rect 1422 538 1427 543
rect 1469 528 1476 535
rect 1569 538 1574 543
rect 1261 511 1266 518
rect 1284 511 1289 518
rect 1407 513 1412 520
rect 1430 513 1435 520
rect 1616 528 1623 535
rect 1554 513 1559 520
rect 1577 513 1582 520
rect 499 427 504 432
rect 605 435 610 441
rect 546 417 553 424
rect 643 427 648 432
rect 745 433 751 440
rect 484 401 489 409
rect 507 402 512 409
rect 690 417 697 424
rect 792 429 797 434
rect 894 436 900 442
rect 839 419 846 426
rect 937 430 942 435
rect 1019 436 1027 443
rect 984 420 991 427
rect 628 402 633 409
rect 651 402 656 409
rect 777 404 782 411
rect 800 404 805 411
rect 922 404 927 411
rect 945 405 950 412
rect 192 357 197 362
rect 272 366 278 371
rect 239 348 246 354
rect 100 326 108 334
rect 177 333 182 340
rect 268 345 277 354
rect 200 334 205 340
rect 17 227 22 232
rect 41 227 47 232
rect 54 227 59 232
rect 77 227 85 232
rect 53 205 59 210
rect 332 347 341 356
rect 191 239 196 244
rect 236 230 244 235
rect 176 214 181 219
rect 198 213 204 219
rect 190 135 195 140
rect 235 126 243 132
rect 190 39 195 44
rect 417 47 427 54
rect 236 29 244 35
rect 198 15 203 22
<< metal2 >>
rect 1240 638 1241 647
rect 591 629 1068 634
rect 591 628 618 629
rect 592 549 598 628
rect 730 621 735 622
rect 730 550 735 614
rect 876 551 881 618
rect 1033 552 1039 599
rect 504 535 530 538
rect 640 535 666 538
rect 786 537 812 540
rect 933 537 959 540
rect 525 531 530 535
rect 525 526 546 531
rect 661 531 666 535
rect 807 533 812 537
rect 661 526 682 531
rect 807 528 828 533
rect 954 533 959 537
rect 954 528 975 533
rect 484 506 489 510
rect 467 501 489 506
rect 507 494 512 510
rect 600 510 620 514
rect 751 512 766 515
rect 751 511 771 512
rect 751 510 767 511
rect 600 509 617 510
rect 643 494 648 510
rect 789 494 794 512
rect 894 515 909 516
rect 894 512 913 515
rect 894 511 918 512
rect 936 494 941 512
rect 1062 506 1068 629
rect 1145 536 1171 539
rect 1166 532 1171 536
rect 1166 527 1187 532
rect 1125 506 1130 511
rect 1062 501 1130 506
rect 1237 515 1241 638
rect 1388 615 1389 624
rect 1281 536 1307 539
rect 1302 532 1307 536
rect 1302 527 1323 532
rect 1236 511 1261 515
rect 1383 517 1389 615
rect 1527 597 1528 604
rect 1427 538 1453 541
rect 1448 534 1453 538
rect 1448 529 1469 534
rect 1383 516 1401 517
rect 1383 513 1407 516
rect 1383 512 1412 513
rect 1523 516 1528 597
rect 1574 538 1600 541
rect 1595 534 1600 538
rect 1595 529 1616 534
rect 422 491 941 494
rect 422 380 426 491
rect 504 427 530 430
rect 525 423 530 427
rect 605 424 610 435
rect 1027 438 1068 443
rect 648 427 674 430
rect 525 418 546 423
rect 669 423 674 427
rect 669 418 690 423
rect 745 412 751 433
rect 797 429 823 432
rect 818 425 823 429
rect 818 420 839 425
rect 896 414 900 436
rect 942 430 968 433
rect 963 426 968 430
rect 963 421 984 426
rect 473 401 484 405
rect 507 380 512 402
rect 618 402 628 405
rect 618 401 633 402
rect 767 404 777 407
rect 767 403 782 404
rect 912 404 922 408
rect 651 380 656 402
rect 800 380 805 404
rect 945 380 950 405
rect 422 377 950 380
rect 278 367 295 371
rect 422 370 426 377
rect 945 376 950 377
rect 418 367 426 370
rect 197 357 223 360
rect 218 353 223 357
rect 218 349 239 353
rect 218 348 230 349
rect 45 326 100 331
rect 177 331 182 333
rect 108 326 182 331
rect 45 234 50 326
rect 200 316 205 334
rect 132 309 205 316
rect 45 232 49 234
rect 132 232 139 309
rect 196 239 219 242
rect 0 227 17 232
rect 47 227 49 232
rect 85 227 139 232
rect 214 235 219 239
rect 223 235 228 348
rect 277 348 332 354
rect 214 230 236 235
rect 0 201 6 227
rect 54 210 58 227
rect 132 215 139 227
rect 132 214 176 215
rect 132 208 181 214
rect 198 201 204 213
rect 0 197 204 201
rect 0 196 6 197
rect 40 15 44 197
rect 195 135 219 138
rect 214 131 219 135
rect 223 131 228 230
rect 214 126 235 131
rect 195 39 218 42
rect 214 35 218 39
rect 223 35 228 126
rect 418 54 422 367
rect 1148 334 1153 511
rect 1284 349 1289 511
rect 1430 365 1435 513
rect 1522 513 1554 516
rect 1522 512 1559 513
rect 1577 495 1582 513
rect 1578 446 1582 495
rect 214 30 236 35
rect 40 12 203 15
rect 198 11 203 12
<< m3contact >>
rect 1033 599 1041 607
rect 1518 597 1527 607
rect 1068 436 1078 444
rect 605 418 610 424
rect 744 405 751 412
rect 895 407 901 414
rect 1577 437 1587 446
rect 1428 357 1438 365
rect 1281 342 1291 349
rect 1148 326 1155 334
<< metal3 >>
rect 1041 605 1051 606
rect 1041 600 1518 605
rect 1041 599 1051 600
rect 1073 444 1577 446
rect 1078 437 1577 444
rect 605 329 610 418
rect 744 349 751 405
rect 895 362 901 407
rect 895 357 1428 362
rect 744 343 1281 349
rect 605 326 1148 329
rect 605 325 1154 326
<< labels >>
rlabel metal1 38 230 38 230 1 S0c
rlabel metal1 23 230 23 230 1 S0
rlabel metal1 61 231 61 231 1 S1
rlabel metal1 277 250 277 250 1 D1
rlabel metal1 271 369 271 369 1 D0
rlabel metal1 279 50 279 50 1 D3
rlabel metal1 188 33 188 33 1 DEC_AND_NODE_4
rlabel metal1 188 56 188 56 1 DEC_D3_NAND
rlabel metal1 280 146 280 146 1 D2
rlabel metal1 189 129 189 129 1 DEC_AND_NODE_3
rlabel metal1 189 152 189 152 1 DEC_D2_NAND
rlabel metal1 191 233 191 233 1 Dec_AND_node_2
rlabel metal1 192 256 192 256 1 DEC_D1_NAND
rlabel metal1 187 375 187 375 1 DEC_D0_NAND
rlabel metal1 192 352 192 352 1 Dec_AND_node_1
rlabel m2contact 80 230 80 230 1 S1c
rlabel metal1 80 212 80 212 1 gnd
rlabel metal1 56 256 56 256 1 vdd
rlabel metal2 479 403 479 403 1 B3
rlabel metal2 620 404 620 404 1 B2
rlabel metal2 772 406 772 406 1 B1
rlabel metal2 915 406 915 406 1 B0
rlabel metal1 938 424 938 424 1 ander_node_5
rlabel metal1 790 424 790 424 1 ander_node_6
rlabel metal1 641 420 641 420 1 ander_node_7
rlabel metal1 496 422 496 422 1 ander_node_8
rlabel metal1 972 441 972 441 1 and_b0e_nand
rlabel metal1 837 440 837 440 1 and_b1e_nand
rlabel metal1 683 437 683 437 1 and_b2e_nand
rlabel metal1 535 437 535 437 1 and_b3e_nand
rlabel metal1 1016 441 1016 441 1 and_b0e
rlabel metal1 872 440 872 440 1 and_b1e
rlabel metal1 724 437 724 437 1 and_b2e
rlabel metal1 580 438 580 438 1 and_b3e
rlabel metal1 1007 547 1007 547 1 and_a0e
rlabel metal1 860 547 860 547 1 and_a1e
rlabel metal1 713 545 713 545 1 and_a2e
rlabel metal1 578 546 578 546 1 and_a3e
rlabel metal1 970 547 970 547 1 and_a0e_nand
rlabel metal1 824 548 824 548 1 and_a1e_nand
rlabel metal1 681 546 681 546 1 and_a2e_nand
rlabel metal1 537 547 537 547 1 and_a3e_nand
rlabel metal1 927 531 927 531 1 ander_node_4
rlabel metal1 780 531 780 531 1 ander_node_3
rlabel metal1 634 530 634 530 1 ander_node_2
rlabel metal1 498 529 498 529 1 ander_node_1
rlabel metal2 907 513 907 513 1 A0
rlabel metal2 761 513 761 513 1 A1
rlabel metal2 614 511 614 511 1 A2
rlabel metal2 486 506 486 506 1 A3
rlabel metal1 1138 531 1138 531 1 ander_node_9
rlabel metal1 1272 531 1272 531 1 ander_node_10
rlabel metal1 1422 534 1422 534 1 ander_node_11
rlabel metal1 1566 531 1566 531 1 ander_node_12
rlabel metal1 1179 547 1179 547 1 A3_and_B3_nand
rlabel metal1 1307 548 1307 548 1 A2_and_B2_nand
rlabel metal1 1462 549 1462 549 1 A1_and_B1_nand
rlabel metal1 1602 549 1602 549 1 A0_and_B0_nand
rlabel metal1 1220 547 1220 547 1 A3_and_B3
rlabel metal1 1356 547 1356 547 1 A2_and_B2
rlabel metal1 1501 549 1501 549 1 A1_and_B1
rlabel metal1 1649 549 1649 549 1 A0_and_B0
<< end >>
