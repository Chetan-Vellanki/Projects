magic
tech scmos
timestamp 1701376110
<< nwell >>
rect -1091 577 -1027 578
rect -1202 558 -1156 577
rect -1131 558 -1027 577
rect 465 566 525 583
rect -1080 551 -1027 558
rect -1079 550 -1027 551
rect 539 550 585 569
rect 600 566 661 583
rect 675 550 721 569
rect 746 568 807 585
rect 821 552 867 571
rect 894 568 954 585
rect 968 552 1014 571
rect 1105 567 1166 584
rect 1180 551 1226 570
rect 1241 567 1302 584
rect 1316 551 1362 570
rect 1387 569 1448 586
rect 1462 553 1508 572
rect 1534 569 1595 586
rect 1609 553 1655 572
rect -1012 511 -945 539
rect -930 515 -884 534
rect 464 458 525 475
rect 539 442 585 461
rect 608 458 669 475
rect 683 442 729 461
rect 757 460 818 477
rect 832 444 878 463
rect 902 461 963 478
rect 977 445 1023 464
rect 157 388 218 405
rect 230 373 276 392
rect -1094 355 -1030 356
rect -1205 336 -1159 355
rect -1134 336 -1030 355
rect -1083 329 -1030 336
rect -710 330 -664 349
rect -650 346 -589 363
rect -563 330 -517 349
rect -503 346 -442 363
rect -1082 328 -1030 329
rect -417 328 -371 347
rect -357 344 -296 361
rect -281 328 -235 347
rect -221 344 -160 361
rect -1008 317 -985 322
rect -1015 289 -948 317
rect -933 293 -887 312
rect 156 270 217 287
rect -719 223 -673 242
rect -659 239 -598 256
rect -574 222 -528 241
rect -514 238 -453 255
rect 229 254 275 273
rect -425 220 -379 239
rect -365 236 -304 253
rect -281 220 -235 239
rect -221 236 -160 253
rect 2 234 86 253
rect -1339 182 -1241 183
rect -1385 163 -1241 182
rect -1091 170 -1027 171
rect -1339 154 -1241 163
rect -1227 151 -1156 170
rect -1131 151 -1027 170
rect 155 166 216 183
rect -1080 144 -1027 151
rect 230 150 276 169
rect -1079 143 -1027 144
rect -1000 135 -982 137
rect -1005 132 -982 135
rect -1012 104 -945 132
rect -930 108 -884 127
rect 155 70 216 87
rect 228 54 275 73
rect -1091 -5 -1027 -4
rect -1202 -24 -1156 -5
rect -1131 -24 -1027 -5
rect -1080 -31 -1027 -24
rect -1079 -32 -1027 -31
rect -1009 -43 -982 -38
rect -1012 -71 -945 -43
rect -930 -67 -884 -48
<< ntransistor >>
rect -982 561 -977 566
rect -964 561 -959 566
rect -1176 543 -1171 548
rect -1116 543 -1111 548
rect 484 543 489 548
rect 507 543 512 548
rect -1065 522 -1060 527
rect -1047 522 -1042 527
rect 620 543 625 548
rect 643 543 648 548
rect 766 545 771 550
rect 789 545 794 550
rect 565 535 570 540
rect 701 535 706 540
rect 913 545 918 550
rect 936 545 941 550
rect 847 537 852 542
rect 1125 544 1130 549
rect 1148 544 1153 549
rect 994 537 999 542
rect 1261 544 1266 549
rect 1284 544 1289 549
rect 1407 546 1412 551
rect 1430 546 1435 551
rect 1206 536 1211 541
rect 1342 536 1347 541
rect 1554 546 1559 551
rect 1577 546 1582 551
rect 1488 538 1493 543
rect 1635 538 1640 543
rect -904 500 -899 505
rect 484 435 489 440
rect 507 435 512 440
rect 628 435 633 440
rect 651 435 656 440
rect 777 437 782 442
rect 800 437 805 442
rect 922 438 927 443
rect 945 438 950 443
rect 565 427 570 432
rect 709 427 714 432
rect 858 429 863 434
rect 1003 430 1008 435
rect 177 365 182 370
rect 200 365 205 370
rect -985 339 -980 344
rect -967 339 -962 344
rect -1179 321 -1174 326
rect -1119 321 -1114 326
rect -1068 300 -1063 305
rect -1050 300 -1045 305
rect -637 323 -632 328
rect -614 323 -609 328
rect -695 315 -690 320
rect -490 323 -485 328
rect -467 323 -462 328
rect 256 358 261 363
rect -548 315 -543 320
rect -344 321 -339 326
rect -321 321 -316 326
rect -402 313 -397 318
rect -208 321 -203 326
rect -185 321 -180 326
rect -266 313 -261 318
rect -907 278 -902 283
rect -646 216 -641 221
rect -623 216 -618 221
rect 176 247 181 252
rect 199 247 204 252
rect -704 208 -699 213
rect -501 215 -496 220
rect -478 215 -473 220
rect 28 219 33 224
rect 66 219 71 224
rect 255 239 260 244
rect -559 207 -554 212
rect -352 213 -347 218
rect -329 213 -324 218
rect -410 205 -405 210
rect -208 213 -203 218
rect -185 213 -180 218
rect -266 205 -261 210
rect -1370 148 -1365 153
rect -982 154 -977 159
rect -964 154 -959 159
rect 175 143 180 148
rect 198 143 203 148
rect -1311 132 -1306 137
rect -1295 132 -1290 137
rect -1279 132 -1274 137
rect -1263 132 -1258 137
rect -1176 136 -1171 141
rect -1116 136 -1111 141
rect -1065 115 -1060 120
rect -1047 115 -1042 120
rect 256 135 261 140
rect -904 93 -899 98
rect 175 47 180 52
rect 198 47 203 52
rect 255 39 260 44
rect -982 -21 -977 -16
rect -964 -21 -959 -16
rect -1176 -39 -1171 -34
rect -1116 -39 -1111 -34
rect -1065 -60 -1060 -55
rect -1047 -60 -1042 -55
rect -904 -82 -899 -77
<< ptransistor >>
rect -1176 565 -1171 570
rect -1116 565 -1111 570
rect 484 572 489 577
rect 507 572 512 577
rect 620 572 625 577
rect 643 572 648 577
rect 766 574 771 579
rect 789 574 794 579
rect 913 574 918 579
rect 936 574 941 579
rect -1065 561 -1060 566
rect -1047 561 -1042 566
rect 565 557 570 562
rect 701 557 706 562
rect 847 559 852 564
rect 1125 573 1130 578
rect 1148 573 1153 578
rect 1261 573 1266 578
rect 1284 573 1289 578
rect 1407 575 1412 580
rect 1430 575 1435 580
rect 1554 575 1559 580
rect 1577 575 1582 580
rect 994 559 999 564
rect -982 522 -977 527
rect -964 522 -959 527
rect -904 522 -899 527
rect 1206 558 1211 563
rect 1342 558 1347 563
rect 1488 560 1493 565
rect 1635 560 1640 565
rect 484 464 489 469
rect 507 464 512 469
rect 628 464 633 469
rect 651 464 656 469
rect 777 466 782 471
rect 800 466 805 471
rect 922 467 927 472
rect 945 467 950 472
rect 565 449 570 454
rect 709 449 714 454
rect 858 451 863 456
rect 1003 452 1008 457
rect 177 394 182 399
rect 200 394 205 399
rect -1179 343 -1174 348
rect -1119 343 -1114 348
rect 256 380 261 385
rect -637 352 -632 357
rect -614 352 -609 357
rect -490 352 -485 357
rect -467 352 -462 357
rect -1068 339 -1063 344
rect -1050 339 -1045 344
rect -695 337 -690 342
rect -548 337 -543 342
rect -344 350 -339 355
rect -321 350 -316 355
rect -208 350 -203 355
rect -185 350 -180 355
rect -402 335 -397 340
rect -985 300 -980 305
rect -967 300 -962 305
rect -907 300 -902 305
rect -266 335 -261 340
rect 176 276 181 281
rect 199 276 204 281
rect -646 245 -641 250
rect -623 245 -618 250
rect -704 230 -699 235
rect -501 244 -496 249
rect -478 244 -473 249
rect 255 261 260 266
rect -559 229 -554 234
rect -352 242 -347 247
rect -329 242 -324 247
rect -208 242 -203 247
rect -185 242 -180 247
rect -410 227 -405 232
rect -266 227 -261 232
rect 28 241 33 246
rect 66 241 71 246
rect -1370 170 -1365 175
rect -1311 166 -1306 171
rect -1295 166 -1290 171
rect -1279 166 -1274 171
rect -1263 166 -1258 171
rect -1176 158 -1171 163
rect -1116 158 -1111 163
rect 175 172 180 177
rect 198 172 203 177
rect -1065 154 -1060 159
rect -1047 154 -1042 159
rect 256 157 261 162
rect -982 115 -977 120
rect -964 115 -959 120
rect -904 115 -899 120
rect 175 76 180 81
rect 198 76 203 81
rect 255 61 260 66
rect -1176 -17 -1171 -12
rect -1116 -17 -1111 -12
rect -1065 -21 -1060 -16
rect -1047 -21 -1042 -16
rect -982 -60 -977 -55
rect -964 -60 -959 -55
rect -904 -60 -899 -55
<< ndiffusion >>
rect -985 561 -982 566
rect -977 561 -964 566
rect -959 561 -956 566
rect -1178 543 -1176 548
rect -1171 543 -1168 548
rect -1119 543 -1116 548
rect -1111 543 -1109 548
rect 482 543 484 548
rect 489 543 491 548
rect 505 543 507 548
rect 512 543 514 548
rect -1068 522 -1065 527
rect -1060 522 -1047 527
rect -1042 522 -1039 527
rect 618 543 620 548
rect 625 543 627 548
rect 641 543 643 548
rect 648 543 650 548
rect 764 545 766 550
rect 771 545 773 550
rect 787 545 789 550
rect 794 545 796 550
rect 563 535 565 540
rect 570 535 573 540
rect 699 535 701 540
rect 706 535 709 540
rect 911 545 913 550
rect 918 545 920 550
rect 934 545 936 550
rect 941 545 943 550
rect 845 537 847 542
rect 852 537 855 542
rect 1123 544 1125 549
rect 1130 544 1132 549
rect 1146 544 1148 549
rect 1153 544 1155 549
rect 992 537 994 542
rect 999 537 1002 542
rect 1259 544 1261 549
rect 1266 544 1268 549
rect 1282 544 1284 549
rect 1289 544 1291 549
rect 1405 546 1407 551
rect 1412 546 1414 551
rect 1428 546 1430 551
rect 1435 546 1437 551
rect 1204 536 1206 541
rect 1211 536 1214 541
rect 1340 536 1342 541
rect 1347 536 1350 541
rect 1552 546 1554 551
rect 1559 546 1561 551
rect 1575 546 1577 551
rect 1582 546 1584 551
rect 1486 538 1488 543
rect 1493 538 1496 543
rect 1633 538 1635 543
rect 1640 538 1643 543
rect -906 500 -904 505
rect -899 500 -896 505
rect 482 435 484 440
rect 489 435 491 440
rect 505 435 507 440
rect 512 435 514 440
rect 626 435 628 440
rect 633 435 635 440
rect 649 435 651 440
rect 656 435 658 440
rect 775 437 777 442
rect 782 437 784 442
rect 798 437 800 442
rect 805 437 807 442
rect 920 438 922 443
rect 927 438 929 443
rect 943 438 945 443
rect 950 438 952 443
rect 563 427 565 432
rect 570 427 573 432
rect 707 427 709 432
rect 714 427 717 432
rect 856 429 858 434
rect 863 429 866 434
rect 1001 430 1003 435
rect 1008 430 1011 435
rect 175 365 177 370
rect 182 365 184 370
rect 198 365 200 370
rect 205 365 207 370
rect -988 339 -985 344
rect -980 339 -967 344
rect -962 339 -959 344
rect -1181 321 -1179 326
rect -1174 321 -1171 326
rect -1122 321 -1119 326
rect -1114 321 -1112 326
rect -1071 300 -1068 305
rect -1063 300 -1050 305
rect -1045 300 -1042 305
rect -639 323 -637 328
rect -632 323 -630 328
rect -616 323 -614 328
rect -609 323 -607 328
rect -698 315 -695 320
rect -690 315 -688 320
rect -492 323 -490 328
rect -485 323 -483 328
rect -469 323 -467 328
rect -462 323 -460 328
rect 254 358 256 363
rect 261 358 264 363
rect -551 315 -548 320
rect -543 315 -541 320
rect -346 321 -344 326
rect -339 321 -337 326
rect -323 321 -321 326
rect -316 321 -314 326
rect -405 313 -402 318
rect -397 313 -395 318
rect -210 321 -208 326
rect -203 321 -201 326
rect -187 321 -185 326
rect -180 321 -178 326
rect -269 313 -266 318
rect -261 313 -259 318
rect -909 278 -907 283
rect -902 278 -899 283
rect -648 216 -646 221
rect -641 216 -639 221
rect -625 216 -623 221
rect -618 216 -616 221
rect 174 247 176 252
rect 181 247 183 252
rect 197 247 199 252
rect 204 247 206 252
rect -707 208 -704 213
rect -699 208 -697 213
rect -503 215 -501 220
rect -496 215 -494 220
rect -480 215 -478 220
rect -473 215 -471 220
rect 26 219 28 224
rect 33 219 36 224
rect 64 219 66 224
rect 71 219 74 224
rect 253 239 255 244
rect 260 239 263 244
rect -562 207 -559 212
rect -554 207 -552 212
rect -354 213 -352 218
rect -347 213 -345 218
rect -331 213 -329 218
rect -324 213 -322 218
rect -413 205 -410 210
rect -405 205 -403 210
rect -210 213 -208 218
rect -203 213 -201 218
rect -187 213 -185 218
rect -180 213 -178 218
rect -269 205 -266 210
rect -261 205 -259 210
rect -1373 148 -1370 153
rect -1365 148 -1363 153
rect -985 154 -982 159
rect -977 154 -964 159
rect -959 154 -956 159
rect 173 143 175 148
rect 180 143 182 148
rect 196 143 198 148
rect 203 143 205 148
rect -1313 132 -1311 137
rect -1306 132 -1295 137
rect -1290 132 -1279 137
rect -1274 132 -1263 137
rect -1258 132 -1255 137
rect -1178 136 -1176 141
rect -1171 136 -1168 141
rect -1119 136 -1116 141
rect -1111 136 -1109 141
rect -1068 115 -1065 120
rect -1060 115 -1047 120
rect -1042 115 -1039 120
rect 254 135 256 140
rect 261 135 264 140
rect -906 93 -904 98
rect -899 93 -896 98
rect 173 47 175 52
rect 180 47 182 52
rect 196 47 198 52
rect 203 47 205 52
rect 253 39 255 44
rect 260 39 263 44
rect -985 -21 -982 -16
rect -977 -21 -964 -16
rect -959 -21 -956 -16
rect -1178 -39 -1176 -34
rect -1171 -39 -1168 -34
rect -1119 -39 -1116 -34
rect -1111 -39 -1109 -34
rect -1068 -60 -1065 -55
rect -1060 -60 -1047 -55
rect -1042 -60 -1039 -55
rect -906 -82 -904 -77
rect -899 -82 -896 -77
<< pdiffusion >>
rect -1178 565 -1176 570
rect -1171 565 -1168 570
rect -1119 565 -1116 570
rect -1111 565 -1109 570
rect 482 572 484 577
rect 489 572 496 577
rect 501 572 507 577
rect 512 572 514 577
rect 618 572 620 577
rect 625 572 632 577
rect 637 572 643 577
rect 648 572 650 577
rect 764 574 766 579
rect 771 574 778 579
rect 783 574 789 579
rect 794 574 796 579
rect 911 574 913 579
rect 918 574 925 579
rect 930 574 936 579
rect 941 574 943 579
rect -1068 561 -1065 566
rect -1060 561 -1047 566
rect -1042 561 -1039 566
rect 563 557 565 562
rect 570 557 573 562
rect 699 557 701 562
rect 706 557 709 562
rect 845 559 847 564
rect 852 559 855 564
rect 1123 573 1125 578
rect 1130 573 1137 578
rect 1142 573 1148 578
rect 1153 573 1155 578
rect 1259 573 1261 578
rect 1266 573 1273 578
rect 1278 573 1284 578
rect 1289 573 1291 578
rect 1405 575 1407 580
rect 1412 575 1419 580
rect 1424 575 1430 580
rect 1435 575 1437 580
rect 1552 575 1554 580
rect 1559 575 1566 580
rect 1571 575 1577 580
rect 1582 575 1584 580
rect 992 559 994 564
rect 999 559 1002 564
rect -985 522 -982 527
rect -977 522 -964 527
rect -959 522 -956 527
rect -906 522 -904 527
rect -899 522 -896 527
rect 1204 558 1206 563
rect 1211 558 1214 563
rect 1340 558 1342 563
rect 1347 558 1350 563
rect 1486 560 1488 565
rect 1493 560 1496 565
rect 1633 560 1635 565
rect 1640 560 1643 565
rect 482 464 484 469
rect 489 464 496 469
rect 501 464 507 469
rect 512 464 514 469
rect 626 464 628 469
rect 633 464 640 469
rect 645 464 651 469
rect 656 464 658 469
rect 775 466 777 471
rect 782 466 789 471
rect 794 466 800 471
rect 805 466 807 471
rect 920 467 922 472
rect 927 467 934 472
rect 939 467 945 472
rect 950 467 952 472
rect 563 449 565 454
rect 570 449 573 454
rect 707 449 709 454
rect 714 449 717 454
rect 856 451 858 456
rect 863 451 866 456
rect 1001 452 1003 457
rect 1008 452 1011 457
rect 175 394 177 399
rect 182 394 189 399
rect 194 394 200 399
rect 205 394 207 399
rect -1181 343 -1179 348
rect -1174 343 -1171 348
rect -1122 343 -1119 348
rect -1114 343 -1112 348
rect 254 380 256 385
rect 261 380 264 385
rect -639 352 -637 357
rect -632 352 -626 357
rect -621 352 -614 357
rect -609 352 -607 357
rect -492 352 -490 357
rect -485 352 -479 357
rect -474 352 -467 357
rect -462 352 -460 357
rect -1071 339 -1068 344
rect -1063 339 -1050 344
rect -1045 339 -1042 344
rect -698 337 -695 342
rect -690 337 -688 342
rect -551 337 -548 342
rect -543 337 -541 342
rect -346 350 -344 355
rect -339 350 -333 355
rect -328 350 -321 355
rect -316 350 -314 355
rect -210 350 -208 355
rect -203 350 -197 355
rect -192 350 -185 355
rect -180 350 -178 355
rect -405 335 -402 340
rect -397 335 -395 340
rect -988 300 -985 305
rect -980 300 -967 305
rect -962 300 -959 305
rect -909 300 -907 305
rect -902 300 -899 305
rect -269 335 -266 340
rect -261 335 -259 340
rect 174 276 176 281
rect 181 276 188 281
rect 193 276 199 281
rect 204 276 206 281
rect -648 245 -646 250
rect -641 245 -635 250
rect -630 245 -623 250
rect -618 245 -616 250
rect -707 230 -704 235
rect -699 230 -697 235
rect -503 244 -501 249
rect -496 244 -490 249
rect -485 244 -478 249
rect -473 244 -471 249
rect 253 261 255 266
rect 260 261 263 266
rect -562 229 -559 234
rect -554 229 -552 234
rect -354 242 -352 247
rect -347 242 -341 247
rect -336 242 -329 247
rect -324 242 -322 247
rect -210 242 -208 247
rect -203 242 -197 247
rect -192 242 -185 247
rect -180 242 -178 247
rect -413 227 -410 232
rect -405 227 -403 232
rect -269 227 -266 232
rect -261 227 -259 232
rect 26 241 28 246
rect 33 241 36 246
rect 64 241 66 246
rect 71 241 74 246
rect -1373 170 -1370 175
rect -1365 170 -1363 175
rect -1314 166 -1311 171
rect -1306 166 -1303 171
rect -1298 166 -1295 171
rect -1290 166 -1287 171
rect -1282 166 -1279 171
rect -1274 166 -1271 171
rect -1266 166 -1263 171
rect -1258 166 -1255 171
rect -1178 158 -1176 163
rect -1171 158 -1168 163
rect -1119 158 -1116 163
rect -1111 158 -1109 163
rect 173 172 175 177
rect 180 172 187 177
rect 192 172 198 177
rect 203 172 205 177
rect -1068 154 -1065 159
rect -1060 154 -1047 159
rect -1042 154 -1039 159
rect 254 157 256 162
rect 261 157 264 162
rect -985 115 -982 120
rect -977 115 -964 120
rect -959 115 -956 120
rect -906 115 -904 120
rect -899 115 -896 120
rect 173 76 175 81
rect 180 76 187 81
rect 192 76 198 81
rect 203 76 205 81
rect 253 61 255 66
rect 260 61 263 66
rect -1178 -17 -1176 -12
rect -1171 -17 -1168 -12
rect -1119 -17 -1116 -12
rect -1111 -17 -1109 -12
rect -1068 -21 -1065 -16
rect -1060 -21 -1047 -16
rect -1042 -21 -1039 -16
rect -985 -60 -982 -55
rect -977 -60 -964 -55
rect -959 -60 -956 -55
rect -906 -60 -904 -55
rect -899 -60 -896 -55
<< ndcontact >>
rect -990 561 -985 566
rect -956 561 -951 566
rect -1183 543 -1178 548
rect -1168 543 -1163 548
rect -1124 543 -1119 548
rect -1109 543 -1104 548
rect 477 543 482 548
rect 491 543 495 548
rect 501 543 505 548
rect 514 543 519 548
rect -1073 522 -1068 527
rect -1039 522 -1034 527
rect 613 543 618 548
rect 627 543 631 548
rect 637 543 641 548
rect 650 543 655 548
rect 759 545 764 550
rect 773 545 777 550
rect 783 545 787 550
rect 796 545 801 550
rect 558 535 563 540
rect 573 535 578 540
rect 694 535 699 540
rect 709 535 714 540
rect 906 545 911 550
rect 920 545 924 550
rect 930 545 934 550
rect 943 545 948 550
rect 840 537 845 542
rect 855 537 860 542
rect 1118 544 1123 549
rect 1132 544 1136 549
rect 1142 544 1146 549
rect 1155 544 1160 549
rect 987 537 992 542
rect 1002 537 1007 542
rect 1254 544 1259 549
rect 1268 544 1272 549
rect 1278 544 1282 549
rect 1291 544 1296 549
rect 1400 546 1405 551
rect 1414 546 1418 551
rect 1424 546 1428 551
rect 1437 546 1442 551
rect 1199 536 1204 541
rect 1214 536 1219 541
rect 1335 536 1340 541
rect 1350 536 1355 541
rect 1547 546 1552 551
rect 1561 546 1565 551
rect 1571 546 1575 551
rect 1584 546 1589 551
rect 1481 538 1486 543
rect 1496 538 1501 543
rect 1628 538 1633 543
rect 1643 538 1648 543
rect -911 500 -906 505
rect -896 500 -891 505
rect 477 435 482 440
rect 491 435 495 440
rect 501 435 505 440
rect 514 435 519 440
rect 621 435 626 440
rect 635 435 639 440
rect 645 435 649 440
rect 658 435 663 440
rect 770 437 775 442
rect 784 437 788 442
rect 794 437 798 442
rect 807 437 812 442
rect 915 438 920 443
rect 929 438 933 443
rect 939 438 943 443
rect 952 438 957 443
rect 558 427 563 432
rect 573 427 578 432
rect 702 427 707 432
rect 717 427 722 432
rect 851 429 856 434
rect 866 429 871 434
rect 996 430 1001 435
rect 1011 430 1016 435
rect 170 365 175 370
rect 184 365 188 370
rect 194 365 198 370
rect 207 365 212 370
rect -993 339 -988 344
rect -959 339 -954 344
rect -1186 321 -1181 326
rect -1171 321 -1166 326
rect -1127 321 -1122 326
rect -1112 321 -1107 326
rect -1076 300 -1071 305
rect -1042 300 -1037 305
rect -644 323 -639 328
rect -630 323 -626 328
rect -620 323 -616 328
rect -607 323 -602 328
rect -703 315 -698 320
rect -688 315 -683 320
rect -497 323 -492 328
rect -483 323 -479 328
rect -473 323 -469 328
rect -460 323 -455 328
rect 249 358 254 363
rect 264 358 269 363
rect -556 315 -551 320
rect -541 315 -536 320
rect -351 321 -346 326
rect -337 321 -333 326
rect -327 321 -323 326
rect -314 321 -309 326
rect -410 313 -405 318
rect -395 313 -390 318
rect -215 321 -210 326
rect -201 321 -197 326
rect -191 321 -187 326
rect -178 321 -173 326
rect -274 313 -269 318
rect -259 313 -254 318
rect -914 278 -909 283
rect -899 278 -894 283
rect -653 216 -648 221
rect -639 216 -635 221
rect -629 216 -625 221
rect -616 216 -611 221
rect 169 247 174 252
rect 183 247 187 252
rect 193 247 197 252
rect 206 247 211 252
rect -712 208 -707 213
rect -697 208 -692 213
rect -508 215 -503 220
rect -494 215 -490 220
rect -484 215 -480 220
rect -471 215 -466 220
rect 21 219 26 224
rect 36 219 41 224
rect 59 219 64 224
rect 74 219 79 224
rect 248 239 253 244
rect 263 239 268 244
rect -567 207 -562 212
rect -552 207 -547 212
rect -359 213 -354 218
rect -345 213 -341 218
rect -335 213 -331 218
rect -322 213 -317 218
rect -418 205 -413 210
rect -403 205 -398 210
rect -215 213 -210 218
rect -201 213 -197 218
rect -191 213 -187 218
rect -178 213 -173 218
rect -274 205 -269 210
rect -259 205 -254 210
rect -1378 148 -1373 153
rect -1363 148 -1358 153
rect -990 154 -985 159
rect -956 154 -951 159
rect 168 143 173 148
rect 182 143 186 148
rect 192 143 196 148
rect 205 143 210 148
rect -1318 132 -1313 137
rect -1255 132 -1250 137
rect -1183 136 -1178 141
rect -1168 136 -1163 141
rect -1124 136 -1119 141
rect -1109 136 -1104 141
rect -1073 115 -1068 120
rect -1039 115 -1034 120
rect 249 135 254 140
rect 264 135 269 140
rect -911 93 -906 98
rect -896 93 -891 98
rect 168 47 173 52
rect 182 47 186 52
rect 192 47 196 52
rect 205 47 210 52
rect 248 39 253 44
rect 263 39 268 44
rect -990 -21 -985 -16
rect -956 -21 -951 -16
rect -1183 -39 -1178 -34
rect -1168 -39 -1163 -34
rect -1124 -39 -1119 -34
rect -1109 -39 -1104 -34
rect -1073 -60 -1068 -55
rect -1039 -60 -1034 -55
rect -911 -82 -906 -77
rect -896 -82 -891 -77
<< pdcontact >>
rect -1183 565 -1178 570
rect -1168 565 -1163 570
rect -1124 565 -1119 570
rect -1109 565 -1104 570
rect 477 572 482 577
rect 496 572 501 577
rect 514 572 519 577
rect 613 572 618 577
rect 632 572 637 577
rect 650 572 655 577
rect 759 574 764 579
rect 778 574 783 579
rect 796 574 801 579
rect 906 574 911 579
rect 925 574 930 579
rect 943 574 948 579
rect -1073 561 -1068 566
rect -1039 561 -1034 566
rect 558 557 563 562
rect 573 557 578 562
rect 694 557 699 562
rect 709 557 714 562
rect 840 559 845 564
rect 855 559 860 564
rect 1118 573 1123 578
rect 1137 573 1142 578
rect 1155 573 1160 578
rect 1254 573 1259 578
rect 1273 573 1278 578
rect 1291 573 1296 578
rect 1400 575 1405 580
rect 1419 575 1424 580
rect 1437 575 1442 580
rect 1547 575 1552 580
rect 1566 575 1571 580
rect 1584 575 1589 580
rect 987 559 992 564
rect 1002 559 1007 564
rect -990 522 -985 527
rect -956 522 -951 527
rect -911 522 -906 527
rect -896 522 -891 527
rect 1199 558 1204 563
rect 1214 558 1219 563
rect 1335 558 1340 563
rect 1350 558 1355 563
rect 1481 560 1486 565
rect 1496 560 1501 565
rect 1628 560 1633 565
rect 1643 560 1648 565
rect 477 464 482 469
rect 496 464 501 469
rect 514 464 519 469
rect 621 464 626 469
rect 640 464 645 469
rect 658 464 663 469
rect 770 466 775 471
rect 789 466 794 471
rect 807 466 812 471
rect 915 467 920 472
rect 934 467 939 472
rect 952 467 957 472
rect 558 449 563 454
rect 573 449 578 454
rect 702 449 707 454
rect 717 449 722 454
rect 851 451 856 456
rect 866 451 871 456
rect 996 452 1001 457
rect 1011 452 1016 457
rect 170 394 175 399
rect 189 394 194 399
rect 207 394 212 399
rect -1186 343 -1181 348
rect -1171 343 -1166 348
rect -1127 343 -1122 348
rect -1112 343 -1107 348
rect 249 380 254 385
rect 264 380 269 385
rect -644 352 -639 357
rect -626 352 -621 357
rect -607 352 -602 357
rect -497 352 -492 357
rect -479 352 -474 357
rect -460 352 -455 357
rect -1076 339 -1071 344
rect -1042 339 -1037 344
rect -703 337 -698 342
rect -688 337 -683 342
rect -556 337 -551 342
rect -541 337 -536 342
rect -351 350 -346 355
rect -333 350 -328 355
rect -314 350 -309 355
rect -215 350 -210 355
rect -197 350 -192 355
rect -178 350 -173 355
rect -410 335 -405 340
rect -395 335 -390 340
rect -993 300 -988 305
rect -959 300 -954 305
rect -914 300 -909 305
rect -899 300 -894 305
rect -274 335 -269 340
rect -259 335 -254 340
rect 169 276 174 281
rect 188 276 193 281
rect 206 276 211 281
rect -653 245 -648 250
rect -635 245 -630 250
rect -616 245 -611 250
rect -712 230 -707 235
rect -697 230 -692 235
rect -508 244 -503 249
rect -490 244 -485 249
rect -471 244 -466 249
rect 248 261 253 266
rect 263 261 268 266
rect -567 229 -562 234
rect -552 229 -547 234
rect -359 242 -354 247
rect -341 242 -336 247
rect -322 242 -317 247
rect -215 242 -210 247
rect -197 242 -192 247
rect -178 242 -173 247
rect -418 227 -413 232
rect -403 227 -398 232
rect -274 227 -269 232
rect -259 227 -254 232
rect 21 241 26 246
rect 36 241 41 246
rect 59 241 64 246
rect 74 241 79 246
rect -1378 170 -1373 175
rect -1363 170 -1358 175
rect -1319 166 -1314 171
rect -1303 166 -1298 171
rect -1287 166 -1282 171
rect -1271 166 -1266 171
rect -1255 166 -1250 171
rect -1183 158 -1178 163
rect -1168 158 -1163 163
rect -1124 158 -1119 163
rect -1109 158 -1104 163
rect 168 172 173 177
rect 187 172 192 177
rect 205 172 210 177
rect -1073 154 -1068 159
rect -1039 154 -1034 159
rect 249 157 254 162
rect 264 157 269 162
rect -990 115 -985 120
rect -956 115 -951 120
rect -911 115 -906 120
rect -896 115 -891 120
rect 168 76 173 81
rect 187 76 192 81
rect 205 76 210 81
rect 248 61 253 66
rect 263 61 268 66
rect -1183 -17 -1178 -12
rect -1168 -17 -1163 -12
rect -1124 -17 -1119 -12
rect -1109 -17 -1104 -12
rect -1073 -21 -1068 -16
rect -1039 -21 -1034 -16
rect -990 -60 -985 -55
rect -956 -60 -951 -55
rect -911 -60 -906 -55
rect -896 -60 -891 -55
<< nsubstratencontact >>
rect -1195 565 -1190 570
rect -1097 565 -1092 570
rect 468 572 473 577
rect 604 572 609 577
rect 751 574 755 579
rect 897 574 902 579
rect -1085 561 -1080 566
rect 546 557 551 562
rect 682 557 687 562
rect 828 559 833 564
rect 1109 573 1114 578
rect 1245 573 1250 578
rect 1391 575 1396 580
rect 1538 575 1543 580
rect 975 559 980 564
rect -1005 520 -999 526
rect -923 522 -918 527
rect 1187 558 1192 563
rect 1323 558 1328 563
rect 1469 560 1474 565
rect 1616 560 1621 565
rect 468 464 473 469
rect 612 464 617 469
rect 761 466 766 471
rect 906 467 911 472
rect 546 449 551 454
rect 690 449 695 454
rect 839 451 844 456
rect 984 452 989 457
rect 161 394 166 399
rect -1198 343 -1193 348
rect -1100 343 -1095 348
rect 237 380 242 385
rect -598 352 -593 357
rect -451 352 -446 357
rect -1088 339 -1083 344
rect -676 337 -671 342
rect -529 337 -524 342
rect -305 350 -300 355
rect -169 350 -164 355
rect -383 335 -378 340
rect -1008 301 -1002 306
rect -926 300 -921 305
rect -247 335 -242 340
rect 160 276 165 281
rect -607 245 -602 250
rect -685 230 -680 235
rect -462 244 -457 249
rect 236 261 241 266
rect -540 229 -535 234
rect -313 242 -308 247
rect -169 242 -164 247
rect -391 227 -386 232
rect -247 227 -242 232
rect 9 241 14 246
rect -1351 170 -1346 175
rect -1331 166 -1326 171
rect -1220 158 -1215 163
rect -1097 158 -1092 163
rect 159 172 164 177
rect -1085 154 -1080 159
rect 237 157 242 162
rect -1005 113 -1000 119
rect -923 115 -918 120
rect 159 76 164 81
rect 236 61 241 66
rect -1195 -17 -1190 -12
rect -1097 -17 -1092 -12
rect -1085 -21 -1080 -16
rect -1005 -60 -1000 -55
rect -923 -60 -918 -55
<< polysilicon >>
rect -1047 587 -1009 588
rect -1004 587 -959 588
rect -1047 583 -959 587
rect -1176 570 -1171 573
rect -1116 570 -1111 573
rect -1065 566 -1060 570
rect -1047 566 -1042 583
rect -982 566 -977 570
rect -964 566 -959 583
rect 484 577 489 591
rect 507 577 512 591
rect 620 577 625 591
rect 643 577 648 591
rect 766 579 771 593
rect 789 579 794 593
rect 913 579 918 593
rect 936 579 941 593
rect 1125 578 1130 592
rect 1148 578 1153 592
rect 1261 578 1266 592
rect 1284 578 1289 592
rect 1407 580 1412 594
rect 1430 580 1435 594
rect 1554 580 1559 594
rect 1577 580 1582 594
rect -1176 556 -1171 565
rect -1175 552 -1171 556
rect -1176 548 -1171 552
rect -1116 556 -1111 565
rect -1116 552 -1112 556
rect -1116 548 -1111 552
rect -1065 549 -1060 561
rect -1047 557 -1042 561
rect -982 549 -977 561
rect -964 557 -959 561
rect -1064 544 -1042 549
rect -982 544 -959 549
rect 484 548 489 572
rect 507 548 512 572
rect 565 562 570 565
rect 565 548 570 557
rect 620 548 625 572
rect 643 548 648 572
rect 701 562 706 565
rect 701 548 706 557
rect 766 550 771 574
rect 789 550 794 574
rect 847 564 852 567
rect 847 550 852 559
rect 913 550 918 574
rect 936 550 941 574
rect 994 564 999 567
rect 994 550 999 559
rect -1176 538 -1171 543
rect -1116 538 -1111 543
rect -1084 532 -1060 537
rect -1084 524 -1079 532
rect -1065 527 -1060 532
rect -1047 527 -1042 544
rect -982 527 -977 531
rect -964 527 -959 544
rect 566 544 570 548
rect -904 527 -899 530
rect -1065 504 -1060 522
rect -1047 516 -1042 522
rect 484 524 489 543
rect -982 504 -977 522
rect -1065 499 -977 504
rect -964 487 -959 522
rect -904 513 -899 522
rect 507 524 512 543
rect 565 540 570 544
rect 702 544 706 548
rect 848 546 852 550
rect 565 530 570 535
rect 620 524 625 543
rect 643 524 648 543
rect 701 540 706 544
rect 701 530 706 535
rect 766 526 771 545
rect 789 526 794 545
rect 847 542 852 546
rect 995 546 999 550
rect 1125 549 1130 573
rect 1148 549 1153 573
rect 1206 563 1211 566
rect 1206 549 1211 558
rect 1261 549 1266 573
rect 1284 549 1289 573
rect 1342 563 1347 566
rect 1342 549 1347 558
rect 1407 551 1412 575
rect 1430 551 1435 575
rect 1488 565 1493 568
rect 1488 551 1493 560
rect 1554 551 1559 575
rect 1577 551 1582 575
rect 1635 565 1640 568
rect 1635 551 1640 560
rect 847 532 852 537
rect 913 526 918 545
rect 936 526 941 545
rect 994 542 999 546
rect 1207 545 1211 549
rect 994 532 999 537
rect 1125 525 1130 544
rect 1148 525 1153 544
rect 1206 541 1211 545
rect 1343 545 1347 549
rect 1489 547 1493 551
rect 1206 531 1211 536
rect 1261 525 1266 544
rect 1284 525 1289 544
rect 1342 541 1347 545
rect 1342 531 1347 536
rect 1407 527 1412 546
rect 1430 527 1435 546
rect 1488 543 1493 547
rect 1636 547 1640 551
rect 1488 533 1493 538
rect 1554 527 1559 546
rect 1577 527 1582 546
rect 1635 543 1640 547
rect 1635 533 1640 538
rect -903 509 -899 513
rect -904 505 -899 509
rect -904 495 -899 500
rect 484 469 489 483
rect 507 469 512 483
rect 628 469 633 483
rect 651 469 656 483
rect 777 471 782 485
rect 800 471 805 485
rect 922 472 927 486
rect 945 472 950 486
rect 484 440 489 464
rect 507 440 512 464
rect 565 454 570 457
rect 565 440 570 449
rect 628 440 633 464
rect 651 440 656 464
rect 709 454 714 457
rect 709 440 714 449
rect 777 442 782 466
rect 800 442 805 466
rect 858 456 863 459
rect 858 442 863 451
rect 922 443 927 467
rect 945 443 950 467
rect 1003 457 1008 460
rect 1003 443 1008 452
rect 566 436 570 440
rect 484 416 489 435
rect 177 399 182 413
rect 200 399 205 413
rect 507 416 512 435
rect 565 432 570 436
rect 710 436 714 440
rect 859 438 863 442
rect 1004 439 1008 443
rect 565 422 570 427
rect 628 416 633 435
rect 651 416 656 435
rect 709 432 714 436
rect 709 422 714 427
rect 777 418 782 437
rect 800 418 805 437
rect 858 434 863 438
rect 858 424 863 429
rect 922 419 927 438
rect 945 419 950 438
rect 1003 435 1008 439
rect 1003 425 1008 430
rect -1050 365 -1012 366
rect -1007 365 -962 366
rect -1050 361 -962 365
rect -1179 348 -1174 351
rect -1119 348 -1114 351
rect -1068 344 -1063 348
rect -1050 344 -1045 361
rect -985 344 -980 348
rect -967 344 -962 361
rect -637 357 -632 371
rect -614 357 -609 371
rect -490 357 -485 371
rect -467 357 -462 371
rect 177 370 182 394
rect 200 370 205 394
rect 256 385 261 388
rect 256 371 261 380
rect -344 355 -339 369
rect -321 355 -316 369
rect -208 355 -203 369
rect -185 355 -180 369
rect 257 367 261 371
rect -1179 334 -1174 343
rect -1178 330 -1174 334
rect -1179 326 -1174 330
rect -1119 334 -1114 343
rect -695 342 -690 345
rect -1119 330 -1115 334
rect -1119 326 -1114 330
rect -1068 327 -1063 339
rect -1050 335 -1045 339
rect -985 327 -980 339
rect -967 335 -962 339
rect -695 328 -690 337
rect -637 328 -632 352
rect -614 328 -609 352
rect -548 342 -543 345
rect -548 328 -543 337
rect -490 328 -485 352
rect -467 328 -462 352
rect -402 340 -397 343
rect -1067 322 -1045 327
rect -985 322 -962 327
rect -1179 316 -1174 321
rect -1119 316 -1114 321
rect -1087 310 -1063 315
rect -1087 302 -1082 310
rect -1068 305 -1063 310
rect -1050 305 -1045 322
rect -985 305 -980 309
rect -967 305 -962 322
rect -695 324 -691 328
rect -695 320 -690 324
rect -548 324 -544 328
rect -695 310 -690 315
rect -907 305 -902 308
rect -637 304 -632 323
rect -1068 282 -1063 300
rect -1050 294 -1045 300
rect -985 282 -980 300
rect -1068 277 -980 282
rect -967 265 -962 300
rect -907 291 -902 300
rect -614 304 -609 323
rect -548 320 -543 324
rect -402 326 -397 335
rect -344 326 -339 350
rect -321 326 -316 350
rect -266 340 -261 343
rect -266 326 -261 335
rect -208 326 -203 350
rect -185 326 -180 350
rect 177 346 182 365
rect 200 346 205 365
rect 256 363 261 367
rect 256 354 261 358
rect -548 310 -543 315
rect -490 304 -485 323
rect -467 304 -462 323
rect -402 322 -398 326
rect -402 318 -397 322
rect -266 322 -262 326
rect -402 308 -397 313
rect -344 302 -339 321
rect -321 302 -316 321
rect -266 318 -261 322
rect -266 308 -261 313
rect -208 302 -203 321
rect -185 302 -180 321
rect -906 287 -902 291
rect -907 283 -902 287
rect 176 281 181 295
rect 199 281 204 295
rect -907 273 -902 278
rect -646 250 -641 264
rect -623 250 -618 264
rect -501 249 -496 263
rect -478 249 -473 263
rect -704 235 -699 238
rect -704 221 -699 230
rect -646 221 -641 245
rect -623 221 -618 245
rect -352 247 -347 261
rect -329 247 -324 261
rect -208 247 -203 261
rect -185 247 -180 261
rect 176 252 181 276
rect 199 252 204 276
rect 255 266 260 269
rect 255 252 260 261
rect -559 234 -554 237
rect -704 217 -700 221
rect -704 213 -699 217
rect -559 220 -554 229
rect -501 220 -496 244
rect -478 220 -473 244
rect 28 246 33 249
rect 66 246 71 249
rect 256 248 260 252
rect -410 232 -405 235
rect -559 216 -555 220
rect -704 203 -699 208
rect -646 197 -641 216
rect -623 197 -618 216
rect -559 212 -554 216
rect -410 218 -405 227
rect -352 218 -347 242
rect -329 218 -324 242
rect -266 232 -261 235
rect -266 218 -261 227
rect -208 218 -203 242
rect -185 218 -180 242
rect 28 232 33 241
rect 66 232 71 241
rect 29 228 33 232
rect 67 228 71 232
rect 28 224 33 228
rect 66 224 71 228
rect 176 228 181 247
rect 199 228 204 247
rect 255 244 260 248
rect 255 234 260 239
rect -559 202 -554 207
rect -501 196 -496 215
rect -478 196 -473 215
rect -410 214 -406 218
rect -410 210 -405 214
rect -266 214 -262 218
rect -410 200 -405 205
rect -352 194 -347 213
rect -1370 175 -1365 178
rect -1311 171 -1306 190
rect -1295 171 -1290 190
rect -329 194 -324 213
rect -266 210 -261 214
rect 28 214 33 219
rect 66 214 71 219
rect -266 200 -261 205
rect -208 194 -203 213
rect -185 194 -180 213
rect -1047 180 -1009 181
rect -1004 180 -959 181
rect -1047 176 -959 180
rect 175 177 180 191
rect 198 177 203 191
rect -1279 171 -1274 175
rect -1263 171 -1258 175
rect -1370 161 -1365 170
rect -1370 157 -1366 161
rect -1370 153 -1365 157
rect -1370 143 -1365 148
rect -1311 137 -1306 166
rect -1295 137 -1290 166
rect -1279 137 -1274 166
rect -1263 137 -1258 166
rect -1176 163 -1171 166
rect -1116 163 -1111 166
rect -1065 159 -1060 163
rect -1047 159 -1042 176
rect -982 159 -977 163
rect -964 159 -959 176
rect -1176 149 -1171 158
rect -1175 145 -1171 149
rect -1176 141 -1171 145
rect -1116 149 -1111 158
rect -1116 145 -1112 149
rect -1116 141 -1111 145
rect -1065 142 -1060 154
rect -1047 150 -1042 154
rect -982 142 -977 154
rect -964 150 -959 154
rect 175 148 180 172
rect 198 148 203 172
rect 256 162 261 165
rect 256 148 261 157
rect 257 144 261 148
rect -1064 137 -1042 142
rect -982 137 -959 142
rect -1311 125 -1306 132
rect -1295 125 -1290 132
rect -1279 115 -1274 132
rect -1263 115 -1258 132
rect -1176 131 -1171 136
rect -1116 131 -1111 136
rect -1084 125 -1060 130
rect -1084 117 -1079 125
rect -1065 120 -1060 125
rect -1047 120 -1042 137
rect -982 120 -977 124
rect -964 120 -959 137
rect 175 124 180 143
rect -904 120 -899 123
rect -1065 97 -1060 115
rect -1047 109 -1042 115
rect 198 124 203 143
rect 256 140 261 144
rect 256 130 261 135
rect -982 97 -977 115
rect -1065 92 -977 97
rect -964 80 -959 115
rect -904 106 -899 115
rect -903 102 -899 106
rect -904 98 -899 102
rect -904 88 -899 93
rect 175 81 180 95
rect 198 81 203 95
rect 175 52 180 76
rect 198 52 203 76
rect 255 66 260 69
rect 255 52 260 61
rect 256 48 260 52
rect 175 28 180 47
rect 198 28 203 47
rect 255 44 260 48
rect 255 34 260 39
rect -1047 5 -1009 6
rect -1004 5 -959 6
rect -1047 1 -959 5
rect -1176 -12 -1171 -9
rect -1116 -12 -1111 -9
rect -1065 -16 -1060 -12
rect -1047 -16 -1042 1
rect -982 -16 -977 -12
rect -964 -16 -959 1
rect -1176 -26 -1171 -17
rect -1175 -30 -1171 -26
rect -1176 -34 -1171 -30
rect -1116 -26 -1111 -17
rect -1116 -30 -1112 -26
rect -1116 -34 -1111 -30
rect -1065 -33 -1060 -21
rect -1047 -25 -1042 -21
rect -982 -33 -977 -21
rect -964 -25 -959 -21
rect -1064 -38 -1042 -33
rect -982 -38 -959 -33
rect -1176 -44 -1171 -39
rect -1116 -44 -1111 -39
rect -1084 -50 -1060 -45
rect -1084 -58 -1079 -50
rect -1065 -55 -1060 -50
rect -1047 -55 -1042 -38
rect -982 -55 -977 -51
rect -964 -55 -959 -38
rect -904 -55 -899 -52
rect -1065 -78 -1060 -60
rect -1047 -66 -1042 -60
rect -982 -78 -977 -60
rect -1065 -83 -977 -78
rect -964 -95 -959 -60
rect -904 -69 -899 -60
rect -903 -73 -899 -69
rect -904 -77 -899 -73
rect -904 -87 -899 -82
<< polycontact >>
rect -1009 587 -1004 592
rect -1180 552 -1175 556
rect -1112 552 -1107 556
rect -1069 544 -1064 549
rect 561 544 566 548
rect -1084 519 -1079 524
rect 484 518 489 524
rect 697 544 702 548
rect 843 546 848 550
rect 507 518 512 524
rect 620 518 625 524
rect 643 518 648 524
rect 766 520 771 526
rect 990 546 995 550
rect 789 520 794 526
rect 913 520 918 526
rect 1202 545 1207 549
rect 936 520 941 526
rect 1125 519 1130 525
rect 1338 545 1343 549
rect 1484 547 1489 551
rect 1148 519 1153 525
rect 1261 519 1266 525
rect 1284 519 1289 525
rect 1407 521 1412 527
rect 1631 547 1636 551
rect 1430 521 1435 527
rect 1554 521 1559 527
rect 1577 521 1582 527
rect -908 509 -903 513
rect -964 482 -959 487
rect 561 436 566 440
rect 484 410 489 416
rect 705 436 710 440
rect 854 438 859 442
rect 999 439 1004 443
rect 507 410 512 416
rect 628 410 633 416
rect 651 410 656 416
rect 777 412 782 418
rect 800 412 805 418
rect 922 413 927 419
rect 945 413 950 419
rect -1012 365 -1007 370
rect 252 367 257 371
rect -1183 330 -1178 334
rect -1115 330 -1110 334
rect -1072 322 -1067 327
rect -1087 297 -1082 302
rect -691 324 -686 328
rect -544 324 -539 328
rect -637 298 -632 304
rect 177 340 182 346
rect 200 340 205 346
rect -614 298 -609 304
rect -490 298 -485 304
rect -398 322 -393 326
rect -262 322 -257 326
rect -467 298 -462 304
rect -344 296 -339 302
rect -321 296 -316 302
rect -208 296 -203 302
rect -185 296 -180 302
rect -911 287 -906 291
rect -967 260 -962 265
rect -700 217 -695 221
rect 251 248 256 252
rect -555 216 -550 220
rect -1311 190 -1305 197
rect -1295 190 -1289 197
rect -646 191 -641 197
rect 24 228 29 232
rect 62 228 67 232
rect 176 222 181 228
rect 199 222 204 228
rect -623 191 -618 197
rect -501 190 -496 196
rect -406 214 -401 218
rect -262 214 -257 218
rect -478 190 -473 196
rect -352 188 -347 194
rect -329 188 -324 194
rect -208 188 -203 194
rect -185 188 -180 194
rect -1009 180 -1004 185
rect -1366 157 -1361 161
rect -1180 145 -1175 149
rect -1112 145 -1107 149
rect 252 144 257 148
rect -1069 137 -1064 142
rect -1279 109 -1272 115
rect -1263 109 -1256 115
rect -1084 112 -1079 117
rect 175 118 180 124
rect 198 118 203 124
rect -908 102 -903 106
rect -964 75 -959 80
rect 251 48 256 52
rect 175 22 180 28
rect 198 22 203 28
rect -1009 5 -1004 10
rect -1180 -30 -1175 -26
rect -1112 -30 -1107 -26
rect -1069 -38 -1064 -33
rect -1084 -63 -1079 -58
rect -908 -73 -903 -69
rect -964 -100 -959 -95
<< metal1 >>
rect -928 607 -927 613
rect -1312 198 -1306 607
rect -711 613 -705 616
rect -913 607 -705 613
rect -1009 594 -872 599
rect -1210 590 -1016 594
rect -1210 556 -1205 590
rect -1195 578 -1032 582
rect -1195 577 -1080 578
rect -1195 570 -1190 577
rect -1183 570 -1178 577
rect -1109 570 -1104 577
rect -1168 556 -1163 565
rect -1097 570 -1092 577
rect -1085 566 -1080 577
rect -1210 553 -1180 556
rect -1184 552 -1180 553
rect -1168 552 -1159 556
rect -1124 556 -1119 565
rect -1073 566 -1068 578
rect -1150 552 -1119 556
rect -1107 552 -1101 556
rect -1168 548 -1163 552
rect -1183 539 -1178 543
rect -1192 534 -1161 539
rect -1150 488 -1146 552
rect -1124 548 -1119 552
rect -1094 552 -1086 556
rect -1090 549 -1086 552
rect -1039 555 -1034 561
rect -1021 555 -1016 590
rect -1009 592 -1004 594
rect -990 572 -937 578
rect -990 566 -985 572
rect -956 555 -951 561
rect -1039 550 -951 555
rect -1090 544 -1069 549
rect -1109 539 -1104 543
rect -1133 534 -1095 539
rect -1105 497 -1100 534
rect -1039 527 -1034 550
rect -1084 516 -1079 519
rect -1005 526 -999 539
rect -1073 497 -1068 522
rect -990 527 -985 537
rect -956 527 -951 550
rect -942 497 -937 572
rect -925 534 -882 539
rect -923 527 -918 534
rect -911 527 -906 534
rect -896 514 -891 522
rect -877 514 -872 594
rect -911 509 -908 513
rect -896 509 -872 514
rect -896 505 -891 509
rect -1105 496 -937 497
rect -911 496 -906 500
rect -1105 492 -858 496
rect -942 491 -858 492
rect -1150 483 -981 488
rect -986 478 -981 483
rect -964 478 -959 482
rect -986 473 -959 478
rect -1311 197 -1306 198
rect -1295 385 -1164 388
rect -1295 197 -1290 385
rect -1012 372 -875 377
rect -1213 368 -1019 372
rect -1213 334 -1208 368
rect -1198 356 -1035 360
rect -1198 355 -1083 356
rect -1198 348 -1193 355
rect -1186 348 -1181 355
rect -1112 348 -1107 355
rect -1171 334 -1166 343
rect -1100 348 -1095 355
rect -1088 344 -1083 355
rect -1213 331 -1183 334
rect -1187 330 -1183 331
rect -1171 330 -1162 334
rect -1127 334 -1122 343
rect -1076 344 -1071 356
rect -1153 330 -1122 334
rect -1110 332 -1089 334
rect -1110 330 -1102 332
rect -1171 326 -1166 330
rect -1186 317 -1181 321
rect -1195 312 -1164 317
rect -1153 266 -1149 330
rect -1127 326 -1122 330
rect -1096 330 -1089 332
rect -1093 327 -1089 330
rect -1042 333 -1037 339
rect -1024 333 -1019 368
rect -1012 370 -1007 372
rect -993 350 -940 356
rect -993 344 -988 350
rect -959 333 -954 339
rect -1042 328 -954 333
rect -1093 322 -1072 327
rect -1112 317 -1107 321
rect -1136 312 -1098 317
rect -1108 275 -1103 312
rect -1042 305 -1037 328
rect -993 322 -990 325
rect -1000 317 -985 322
rect -1087 294 -1082 297
rect -1008 306 -1003 317
rect -993 305 -988 317
rect -959 305 -954 328
rect -1076 275 -1071 300
rect -945 275 -940 350
rect -928 312 -885 317
rect -926 305 -921 312
rect -914 305 -909 312
rect -899 292 -894 300
rect -880 292 -875 372
rect -914 287 -911 291
rect -899 287 -875 292
rect -865 309 -859 491
rect -818 440 -811 491
rect -768 467 -767 474
rect -768 410 -761 467
rect -836 402 -760 410
rect -711 402 -705 607
rect 288 611 603 615
rect 467 610 603 611
rect 683 608 688 651
rect 730 641 1230 646
rect 730 621 736 641
rect 683 604 744 608
rect 800 607 805 622
rect 883 618 1378 624
rect 800 604 893 607
rect 305 588 312 593
rect 1439 591 1539 592
rect 1586 591 1617 592
rect 798 590 898 591
rect 945 590 976 591
rect 1391 590 1617 591
rect 744 589 976 590
rect 1157 589 1188 590
rect 1293 589 1617 590
rect 516 588 547 589
rect 652 588 976 589
rect 1102 588 1617 589
rect 305 587 1442 588
rect 305 585 801 587
rect 305 583 519 585
rect -649 461 -640 486
rect -649 455 -279 461
rect -599 423 -573 429
rect -286 421 -279 455
rect -661 406 -430 410
rect 83 410 88 412
rect 305 411 312 583
rect 447 582 474 583
rect 447 482 455 582
rect 468 577 473 582
rect 477 577 482 583
rect 514 577 519 583
rect 539 584 655 585
rect 539 574 543 584
rect 604 583 655 584
rect 604 577 609 583
rect 496 562 501 572
rect 539 569 587 574
rect 613 577 618 583
rect 650 577 655 583
rect 675 574 679 585
rect 751 579 755 585
rect 759 579 764 585
rect 796 579 801 585
rect 821 576 825 587
rect 897 585 948 587
rect 897 579 902 585
rect 491 558 501 562
rect 546 562 551 569
rect 491 554 495 558
rect 558 562 563 569
rect 632 562 637 572
rect 675 569 723 574
rect 491 551 532 554
rect 491 548 495 551
rect 529 548 532 551
rect 573 548 578 557
rect 627 558 637 562
rect 682 562 687 569
rect 627 554 631 558
rect 694 562 699 569
rect 778 564 783 574
rect 821 571 869 576
rect 906 579 911 585
rect 943 579 948 585
rect 968 586 1442 587
rect 968 584 1160 586
rect 968 576 972 584
rect 1102 583 1115 584
rect 1109 578 1114 583
rect 627 551 668 554
rect 474 532 477 546
rect 519 543 521 546
rect 529 544 561 548
rect 573 544 592 548
rect 501 540 504 543
rect 518 532 521 543
rect 573 540 578 544
rect 627 548 631 551
rect 665 548 668 551
rect 709 548 714 557
rect 773 560 783 564
rect 828 564 833 571
rect 773 556 777 560
rect 840 564 845 571
rect 925 564 930 574
rect 968 571 1016 576
rect 1118 578 1123 584
rect 1155 578 1160 584
rect 1180 585 1296 586
rect 1180 575 1184 585
rect 1245 584 1296 585
rect 1245 578 1250 584
rect 773 553 814 556
rect 773 550 777 553
rect 811 550 814 553
rect 855 550 860 559
rect 920 560 930 564
rect 975 564 980 571
rect 920 556 924 560
rect 987 564 992 571
rect 1137 563 1142 573
rect 1180 570 1228 575
rect 1254 578 1259 584
rect 1291 578 1296 584
rect 1316 575 1320 586
rect 1391 580 1396 586
rect 1400 580 1405 586
rect 1437 580 1442 586
rect 1462 577 1466 588
rect 1538 586 1589 588
rect 1538 580 1543 586
rect 920 553 961 556
rect 474 527 521 532
rect 558 531 563 535
rect 610 532 613 546
rect 655 543 657 546
rect 665 544 697 548
rect 709 544 730 548
rect 637 540 640 543
rect 654 532 657 543
rect 709 540 714 544
rect 553 526 588 531
rect 610 527 657 532
rect 484 517 489 518
rect 507 517 512 518
rect 584 505 588 526
rect 694 531 699 535
rect 756 534 759 548
rect 801 545 803 548
rect 811 546 843 550
rect 855 546 876 550
rect 783 542 786 545
rect 800 534 803 545
rect 855 542 860 546
rect 920 550 924 553
rect 958 550 961 553
rect 1002 550 1007 559
rect 1132 559 1142 563
rect 1187 563 1192 570
rect 1132 555 1136 559
rect 1199 563 1204 570
rect 1273 563 1278 573
rect 1316 570 1364 575
rect 1132 552 1173 555
rect 689 530 724 531
rect 689 526 737 530
rect 756 529 803 534
rect 840 533 845 537
rect 903 534 906 548
rect 948 545 950 548
rect 958 546 990 550
rect 1002 546 1032 550
rect 930 542 933 545
rect 947 534 950 545
rect 1002 542 1007 546
rect 1132 549 1136 552
rect 1170 549 1173 552
rect 1214 549 1219 558
rect 1268 559 1278 563
rect 1323 563 1328 570
rect 1268 555 1272 559
rect 1335 563 1340 570
rect 1419 565 1424 575
rect 1462 572 1510 577
rect 1547 580 1552 586
rect 1584 580 1589 586
rect 1609 577 1613 588
rect 1268 552 1309 555
rect 1268 549 1272 552
rect 1306 549 1309 552
rect 1350 549 1355 558
rect 1414 561 1424 565
rect 1469 565 1474 572
rect 1414 557 1418 561
rect 1481 565 1486 572
rect 1566 565 1571 575
rect 1609 572 1657 577
rect 1414 554 1455 557
rect 1414 551 1418 554
rect 1452 551 1455 554
rect 1496 551 1501 560
rect 1561 561 1571 565
rect 1616 565 1621 572
rect 1561 557 1565 561
rect 1628 565 1633 572
rect 1561 554 1602 557
rect 1561 551 1565 554
rect 1599 551 1602 554
rect 1643 551 1648 560
rect 835 528 873 533
rect 903 529 950 534
rect 718 525 737 526
rect 620 517 625 518
rect 643 517 648 518
rect 728 505 735 525
rect 766 519 771 520
rect 789 519 794 520
rect 864 505 873 528
rect 987 533 992 537
rect 1115 533 1118 547
rect 1160 544 1162 547
rect 1170 545 1202 549
rect 1214 545 1222 549
rect 1142 541 1145 544
rect 1159 533 1162 544
rect 1214 541 1219 545
rect 982 528 1018 533
rect 1115 528 1162 533
rect 913 519 918 520
rect 936 519 941 520
rect 1009 505 1018 528
rect 1199 532 1204 536
rect 1251 533 1254 547
rect 1296 544 1298 547
rect 1306 545 1338 549
rect 1350 545 1358 549
rect 1278 541 1281 544
rect 1295 533 1298 544
rect 1350 541 1355 545
rect 1194 527 1229 532
rect 1251 528 1298 533
rect 1125 518 1130 519
rect 1148 518 1153 519
rect 1225 506 1229 527
rect 1335 532 1340 536
rect 1397 535 1400 549
rect 1442 546 1444 549
rect 1452 547 1484 551
rect 1496 547 1504 551
rect 1424 543 1427 546
rect 1441 535 1444 546
rect 1496 543 1501 547
rect 1330 531 1365 532
rect 1330 527 1378 531
rect 1397 530 1444 535
rect 1481 534 1486 538
rect 1544 535 1547 549
rect 1589 546 1591 549
rect 1599 547 1631 551
rect 1643 547 1651 551
rect 1571 543 1574 546
rect 1588 535 1591 546
rect 1643 543 1648 547
rect 1476 529 1514 534
rect 1544 530 1591 535
rect 1359 526 1378 527
rect 1261 518 1266 519
rect 1284 518 1289 519
rect 1369 506 1376 526
rect 1407 520 1412 521
rect 1430 520 1435 521
rect 1505 506 1514 529
rect 1628 534 1633 538
rect 1623 529 1659 534
rect 1554 520 1559 521
rect 1577 520 1582 521
rect 1650 506 1659 529
rect 1037 505 1045 506
rect 584 499 1045 505
rect 1225 501 1660 506
rect 1225 500 1635 501
rect 1037 488 1045 499
rect 1246 488 1255 500
rect 954 483 985 484
rect 809 482 985 483
rect 447 480 477 482
rect 685 481 985 482
rect 516 480 547 481
rect 660 480 985 481
rect 1036 480 1255 488
rect 447 479 957 480
rect 447 477 812 479
rect 821 478 957 479
rect 447 475 519 477
rect 538 475 663 477
rect 468 469 473 475
rect 477 469 482 475
rect 514 469 519 475
rect 539 466 543 475
rect 612 469 617 475
rect 496 454 501 464
rect 539 461 587 466
rect 621 469 626 475
rect 658 469 663 475
rect 683 466 687 477
rect 761 471 766 477
rect 770 471 775 477
rect 807 471 812 477
rect 832 468 836 478
rect 906 472 911 478
rect 491 450 501 454
rect 546 454 551 461
rect 491 446 495 450
rect 558 454 563 461
rect 640 454 645 464
rect 683 461 731 466
rect 491 443 532 446
rect 491 440 495 443
rect 529 440 532 443
rect 573 440 578 449
rect 635 450 645 454
rect 690 454 695 461
rect 635 446 639 450
rect 702 454 707 461
rect 789 456 794 466
rect 832 463 880 468
rect 915 472 920 478
rect 952 472 957 478
rect 977 469 981 480
rect 635 443 676 446
rect 474 424 477 438
rect 519 435 521 438
rect 529 436 561 440
rect 573 436 605 440
rect 501 432 504 435
rect 518 424 521 435
rect 573 432 578 436
rect 635 440 639 443
rect 673 440 676 443
rect 717 440 722 449
rect 784 452 794 456
rect 839 456 844 463
rect 784 448 788 452
rect 851 456 856 463
rect 934 457 939 467
rect 977 464 1025 469
rect 784 445 825 448
rect 784 442 788 445
rect 822 442 825 445
rect 866 442 871 451
rect 929 453 939 457
rect 984 457 989 464
rect 929 449 933 453
rect 996 457 1001 464
rect 929 446 970 449
rect 929 443 933 446
rect 967 443 970 446
rect 1011 443 1016 452
rect 474 419 521 424
rect 558 423 563 427
rect 618 424 621 438
rect 663 435 665 438
rect 673 436 705 440
rect 717 436 745 440
rect 645 432 648 435
rect 662 424 665 435
rect 717 432 722 436
rect 553 418 588 423
rect 618 419 665 424
rect 209 410 312 411
rect 83 407 313 410
rect 83 406 212 407
rect -712 397 -705 402
rect -803 376 -737 383
rect -711 354 -705 397
rect -672 368 -641 369
rect -594 368 -494 369
rect -672 367 -446 368
rect -672 366 -348 367
rect -243 366 -212 367
rect 83 366 88 406
rect 161 405 212 406
rect 161 399 166 405
rect 170 399 175 405
rect 207 399 212 405
rect 232 397 236 407
rect 305 397 313 407
rect 484 409 489 410
rect 507 409 512 410
rect 189 384 194 394
rect 230 392 313 397
rect 184 380 194 384
rect 237 385 242 392
rect 249 385 254 392
rect 184 376 188 380
rect 184 373 225 376
rect 184 370 188 373
rect 222 370 225 373
rect 264 371 269 380
rect 305 372 313 392
rect 229 370 252 371
rect -672 365 88 366
rect -668 354 -664 365
rect -712 349 -664 354
rect -644 363 -593 365
rect -644 357 -639 363
rect -607 357 -602 363
rect -598 357 -593 363
rect -521 354 -517 365
rect -688 342 -683 349
rect -676 342 -671 349
rect -626 342 -621 352
rect -565 349 -517 354
rect -497 363 88 365
rect -497 357 -492 363
rect -460 357 -455 363
rect -451 357 -446 363
rect -375 352 -371 363
rect -541 342 -536 349
rect -626 338 -616 342
rect -703 328 -698 337
rect -620 334 -616 338
rect -657 331 -616 334
rect -657 328 -654 331
rect -620 328 -616 331
rect -529 342 -524 349
rect -479 342 -474 352
rect -419 347 -371 352
rect -351 362 -235 363
rect -351 361 -300 362
rect -351 355 -346 361
rect -314 355 -309 361
rect -305 355 -300 361
rect -239 352 -235 362
rect -479 338 -469 342
rect -395 340 -390 347
rect -721 324 -698 328
rect -686 324 -654 328
rect -703 320 -698 324
rect -646 323 -644 326
rect -688 311 -683 315
rect -646 312 -643 323
rect -629 320 -626 323
rect -602 312 -599 326
rect -556 328 -551 337
rect -473 334 -469 338
rect -510 331 -469 334
rect -510 328 -507 331
rect -473 328 -469 331
rect -383 340 -378 347
rect -333 340 -328 350
rect -283 347 -235 352
rect -215 361 88 363
rect -215 355 -210 361
rect -178 355 -173 361
rect -170 360 88 361
rect -169 355 -164 360
rect -259 340 -254 347
rect -333 336 -323 340
rect -567 325 -551 328
rect -569 324 -551 325
rect -539 324 -507 328
rect -556 320 -551 324
rect -499 323 -497 326
rect -714 309 -678 311
rect -865 306 -678 309
rect -865 304 -705 306
rect -646 307 -599 312
rect -541 311 -536 315
rect -499 312 -496 323
rect -482 320 -479 323
rect -455 312 -452 326
rect -410 326 -405 335
rect -327 332 -323 336
rect -364 329 -323 332
rect -364 326 -361 329
rect -327 326 -323 329
rect -247 340 -242 347
rect -197 340 -192 350
rect -197 336 -187 340
rect -274 326 -269 335
rect -191 332 -187 336
rect -228 329 -187 332
rect -228 326 -225 329
rect -191 326 -187 329
rect -422 322 -405 326
rect -393 322 -361 326
rect -410 318 -405 322
rect -353 321 -351 324
rect -284 325 -269 326
rect -569 306 -531 311
rect -899 283 -894 287
rect -1108 274 -940 275
rect -914 274 -909 278
rect -865 274 -859 304
rect -1108 270 -859 274
rect -945 269 -859 270
rect -1153 261 -984 266
rect -989 256 -984 261
rect -967 256 -962 260
rect -989 251 -962 256
rect -1244 187 -1239 192
rect -1009 187 -872 192
rect -1387 183 -1239 187
rect -1235 183 -1016 187
rect -1387 182 -1339 183
rect -1363 175 -1358 182
rect -1351 175 -1346 182
rect -1331 171 -1326 183
rect -1378 161 -1373 170
rect -1319 171 -1314 183
rect -1287 171 -1282 183
rect -1255 171 -1250 183
rect -1303 163 -1298 166
rect -1318 162 -1298 163
rect -1271 162 -1266 166
rect -1385 157 -1373 161
rect -1361 157 -1342 161
rect -1378 153 -1373 157
rect -1363 144 -1358 148
rect -1346 149 -1342 157
rect -1318 158 -1266 162
rect -1318 149 -1313 158
rect -1346 144 -1313 149
rect -1235 149 -1230 183
rect -1220 171 -1032 175
rect -1220 170 -1080 171
rect -1220 163 -1215 170
rect -1183 163 -1178 170
rect -1109 163 -1104 170
rect -1168 149 -1163 158
rect -1097 163 -1092 170
rect -1085 159 -1080 170
rect -1124 149 -1119 158
rect -1073 159 -1068 171
rect -1235 146 -1180 149
rect -1184 145 -1180 146
rect -1168 145 -1160 149
rect -1388 139 -1349 144
rect -1354 123 -1349 139
rect -1318 137 -1313 144
rect -1168 141 -1163 145
rect -1150 145 -1119 149
rect -1107 147 -1086 149
rect -1107 145 -1100 147
rect -1183 132 -1178 136
rect -1255 130 -1250 132
rect -1217 130 -1161 132
rect -1255 127 -1161 130
rect -1255 126 -1213 127
rect -1255 123 -1250 126
rect -1354 119 -1250 123
rect -1235 112 -1202 115
rect -1279 93 -1274 109
rect -1263 104 -1258 109
rect -1263 100 -1162 104
rect -1279 89 -1245 93
rect -1150 81 -1146 145
rect -1124 141 -1119 145
rect -1095 145 -1086 147
rect -1090 142 -1086 145
rect -1039 148 -1034 154
rect -1021 148 -1016 183
rect -1009 185 -1004 187
rect -990 165 -937 171
rect -990 159 -985 165
rect -956 148 -951 154
rect -1039 143 -951 148
rect -1090 137 -1069 142
rect -1109 132 -1104 136
rect -1133 127 -1095 132
rect -1105 90 -1100 127
rect -1039 120 -1034 143
rect -990 137 -987 140
rect -1084 109 -1079 112
rect -997 132 -982 137
rect -1005 119 -1000 132
rect -1073 90 -1068 115
rect -990 120 -985 132
rect -956 120 -951 143
rect -942 90 -937 165
rect -925 127 -882 132
rect -923 120 -918 127
rect -911 120 -906 127
rect -896 107 -891 115
rect -877 107 -872 187
rect -911 102 -908 106
rect -896 102 -872 107
rect -896 98 -891 102
rect -1105 89 -937 90
rect -911 89 -906 93
rect -865 89 -859 269
rect -847 276 -846 285
rect -741 283 -733 284
rect -714 283 -705 304
rect -637 297 -632 298
rect -614 297 -609 298
rect -569 283 -560 306
rect -499 307 -452 312
rect -395 309 -390 313
rect -353 310 -350 321
rect -336 318 -333 321
rect -309 310 -306 324
rect -279 322 -269 325
rect -257 322 -225 326
rect -274 318 -269 322
rect -217 321 -215 324
rect -420 308 -385 309
rect -433 304 -385 308
rect -490 297 -485 298
rect -433 303 -414 304
rect -353 305 -306 310
rect -259 309 -254 313
rect -217 310 -214 321
rect -200 318 -197 321
rect -173 310 -170 324
rect -284 304 -249 309
rect -467 297 -462 298
rect -431 283 -424 303
rect -344 295 -339 296
rect -321 295 -316 296
rect -284 283 -280 304
rect -217 305 -170 310
rect -208 295 -203 296
rect -185 295 -180 296
rect -847 233 -840 276
rect -813 199 -807 282
rect -741 277 -280 283
rect -843 193 -807 199
rect -770 168 -768 177
rect -770 100 -761 168
rect -1105 85 -857 89
rect -942 84 -857 85
rect -1150 76 -981 81
rect -986 71 -981 76
rect -964 71 -959 75
rect -986 66 -959 71
rect -886 47 -882 69
rect -1009 12 -872 17
rect -1210 8 -1016 12
rect -1210 -26 -1205 8
rect -1195 -4 -1032 0
rect -1195 -5 -1080 -4
rect -1195 -12 -1190 -5
rect -1183 -12 -1178 -5
rect -1109 -12 -1104 -5
rect -1168 -26 -1163 -17
rect -1097 -12 -1092 -5
rect -1085 -16 -1080 -5
rect -1124 -26 -1119 -17
rect -1073 -16 -1068 -4
rect -1210 -29 -1180 -26
rect -1184 -30 -1180 -29
rect -1168 -30 -1160 -26
rect -1168 -34 -1163 -30
rect -1150 -30 -1119 -26
rect -1107 -28 -1086 -26
rect -1107 -30 -1100 -28
rect -1183 -43 -1178 -39
rect -1192 -48 -1161 -43
rect -1150 -94 -1146 -30
rect -1124 -34 -1119 -30
rect -1094 -30 -1086 -28
rect -1090 -33 -1086 -30
rect -1039 -27 -1034 -21
rect -1021 -27 -1016 8
rect -1009 10 -1004 12
rect -990 -10 -937 -4
rect -990 -16 -985 -10
rect -956 -27 -951 -21
rect -1039 -32 -951 -27
rect -1090 -38 -1069 -33
rect -1109 -43 -1104 -39
rect -1133 -48 -1095 -43
rect -1105 -85 -1100 -48
rect -1039 -55 -1034 -32
rect -990 -38 -987 -35
rect -1000 -43 -982 -38
rect -1084 -66 -1079 -63
rect -1009 -55 -1002 -43
rect -990 -55 -985 -43
rect -1009 -60 -1005 -55
rect -956 -55 -951 -32
rect -1073 -85 -1068 -60
rect -942 -85 -937 -10
rect -925 -48 -882 -43
rect -923 -55 -918 -48
rect -911 -55 -906 -48
rect -896 -68 -891 -60
rect -877 -68 -872 12
rect -911 -73 -908 -69
rect -896 -73 -872 -68
rect -896 -77 -891 -73
rect -1105 -86 -937 -85
rect -911 -86 -906 -82
rect -865 -86 -859 84
rect -771 16 -761 100
rect -771 -49 -762 16
rect -1105 -90 -859 -86
rect -942 -91 -859 -90
rect -1150 -99 -981 -94
rect -986 -104 -981 -99
rect -964 -104 -959 -100
rect -986 -109 -959 -104
rect -912 -127 -905 -118
rect -753 -127 -747 217
rect -741 171 -733 277
rect -681 261 -650 262
rect -681 260 -505 261
rect -151 260 -143 360
rect -681 259 -381 260
rect -681 258 -356 259
rect -243 258 -212 259
rect -173 258 -143 260
rect 83 258 88 360
rect 167 354 170 368
rect 212 365 214 368
rect 222 367 252 370
rect 264 367 272 371
rect 222 366 249 367
rect 194 362 197 365
rect 211 354 214 365
rect 264 363 269 367
rect 306 367 312 372
rect 446 367 449 397
rect 580 394 589 418
rect 702 423 707 427
rect 767 426 770 440
rect 812 437 814 440
rect 822 438 854 442
rect 866 438 894 442
rect 794 434 797 437
rect 811 426 814 437
rect 866 434 871 438
rect 697 418 738 423
rect 767 421 814 426
rect 851 425 856 429
rect 912 427 915 441
rect 957 438 959 441
rect 967 439 999 443
rect 1011 439 1019 443
rect 939 435 942 438
rect 956 427 959 438
rect 1011 435 1016 439
rect 846 420 881 425
rect 912 422 959 427
rect 996 426 1001 430
rect 1020 426 1027 427
rect 991 421 1027 426
rect 628 409 633 410
rect 651 409 656 410
rect 730 394 737 418
rect 777 411 782 412
rect 800 411 805 412
rect 874 394 881 420
rect 922 411 927 413
rect 945 412 950 413
rect 1020 394 1027 421
rect 580 393 1027 394
rect 1037 393 1045 480
rect 1246 479 1255 480
rect 580 388 1045 393
rect 249 354 254 358
rect 167 349 214 354
rect 246 349 268 354
rect 261 348 268 349
rect -677 247 -673 258
rect -721 242 -673 247
rect -653 257 -143 258
rect -653 256 -517 257
rect -653 250 -648 256
rect -616 250 -611 256
rect -607 250 -602 256
rect -532 246 -528 256
rect -697 235 -692 242
rect -685 235 -680 242
rect -635 235 -630 245
rect -576 241 -528 246
rect -508 255 -143 257
rect -508 249 -503 255
rect -471 249 -466 255
rect -462 249 -457 255
rect -383 244 -379 255
rect -635 231 -625 235
rect -552 234 -547 241
rect -712 221 -707 230
rect -629 227 -625 231
rect -666 224 -625 227
rect -666 221 -663 224
rect -629 221 -625 224
rect -540 234 -535 241
rect -490 234 -485 244
rect -427 239 -379 244
rect -359 253 -234 255
rect -215 253 -143 255
rect 2 253 88 258
rect 305 353 313 367
rect 304 348 314 353
rect -359 247 -354 253
rect -322 247 -317 253
rect -313 247 -308 253
rect -239 244 -235 253
rect -490 230 -480 234
rect -403 232 -398 239
rect -720 217 -707 221
rect -695 217 -663 221
rect -712 213 -707 217
rect -655 216 -653 219
rect -723 204 -716 205
rect -697 204 -692 208
rect -655 205 -652 216
rect -638 213 -635 216
rect -611 205 -608 219
rect -567 220 -562 229
rect -484 226 -480 230
rect -521 223 -480 226
rect -521 220 -518 223
rect -484 220 -480 223
rect -391 232 -386 239
rect -341 232 -336 242
rect -283 239 -235 244
rect -215 247 -210 253
rect -178 247 -173 253
rect -169 247 -164 253
rect 9 246 14 253
rect -259 232 -254 239
rect -341 228 -331 232
rect -579 217 -562 220
rect -570 216 -562 217
rect -550 216 -518 220
rect -567 212 -562 216
rect -510 215 -508 218
rect -418 218 -413 227
rect -335 224 -331 228
rect -372 221 -331 224
rect -372 218 -369 221
rect -335 218 -331 221
rect -247 232 -242 239
rect -197 232 -192 242
rect 21 246 26 253
rect 59 246 64 253
rect -197 228 -187 232
rect -723 199 -687 204
rect -723 172 -716 199
rect -655 200 -608 205
rect -552 203 -547 207
rect -510 204 -507 215
rect -493 212 -490 215
rect -466 204 -463 218
rect -436 213 -413 218
rect -401 214 -369 218
rect -418 210 -413 213
rect -361 213 -359 216
rect -577 198 -542 203
rect -646 190 -641 191
rect -623 189 -618 191
rect -577 172 -570 198
rect -510 199 -463 204
rect -403 201 -398 205
rect -361 202 -358 213
rect -344 210 -341 213
rect -317 202 -314 216
rect -274 218 -269 227
rect -191 224 -187 228
rect 22 228 24 232
rect 22 227 23 228
rect 36 224 41 241
rect 74 232 79 241
rect 59 228 62 232
rect 74 227 77 232
rect 74 224 79 227
rect -228 221 -187 224
rect -228 218 -225 221
rect -191 218 -187 221
rect -293 214 -269 218
rect -257 214 -225 218
rect -274 210 -269 214
rect -217 213 -215 216
rect -434 196 -393 201
rect -501 189 -496 190
rect -478 189 -473 190
rect -433 172 -426 196
rect -361 197 -314 202
rect -259 201 -254 205
rect -217 202 -214 213
rect -200 210 -197 213
rect -173 202 -170 216
rect 21 215 26 219
rect 59 217 64 219
rect 46 215 65 217
rect -284 196 -249 201
rect -352 187 -347 188
rect -329 187 -324 188
rect -285 172 -276 196
rect -217 197 -170 202
rect 10 214 91 215
rect 10 210 49 214
rect 62 212 91 214
rect 64 210 91 212
rect -208 187 -203 188
rect -185 187 -180 188
rect -139 179 -70 183
rect -723 171 -276 172
rect -741 166 -276 171
rect -723 165 -716 166
rect -433 164 -426 166
rect -285 147 -277 166
rect 10 147 16 210
rect -285 143 17 147
rect -69 -25 -65 15
rect 10 5 16 143
rect 54 106 58 205
rect 100 118 108 326
rect 208 292 239 293
rect 160 289 239 292
rect 160 287 211 289
rect 160 281 165 287
rect 169 281 174 287
rect 206 281 211 287
rect 231 278 235 289
rect 305 278 313 348
rect 547 353 556 355
rect 341 348 556 353
rect 547 319 556 348
rect 688 319 695 388
rect 730 386 737 388
rect 1020 387 1027 388
rect 547 313 696 319
rect 688 311 695 313
rect 188 266 193 276
rect 229 273 313 278
rect 183 262 193 266
rect 236 266 241 273
rect 183 258 187 262
rect 248 266 253 273
rect 286 272 300 273
rect 183 255 224 258
rect 183 252 187 255
rect 221 252 224 255
rect 263 252 268 261
rect 166 236 169 250
rect 211 247 213 250
rect 221 248 251 252
rect 263 248 280 252
rect 193 244 196 247
rect 210 236 213 247
rect 263 244 268 248
rect 166 231 213 236
rect 248 235 253 239
rect 244 230 274 235
rect 176 219 181 222
rect 198 219 204 222
rect 207 188 238 189
rect 159 185 238 188
rect 159 183 210 185
rect 159 177 164 183
rect 168 177 173 183
rect 205 177 210 183
rect 230 174 234 185
rect 305 174 313 273
rect 187 162 192 172
rect 230 169 313 174
rect 182 158 192 162
rect 237 162 242 169
rect 182 154 186 158
rect 249 162 254 169
rect 182 151 223 154
rect 182 148 186 151
rect 220 148 223 151
rect 264 148 269 157
rect 165 132 168 146
rect 210 143 212 146
rect 220 144 252 148
rect 264 144 282 148
rect 192 140 195 143
rect 209 132 212 143
rect 264 140 269 144
rect 165 127 212 132
rect 249 131 254 135
rect 243 126 270 131
rect 100 113 180 118
rect 198 106 203 118
rect 54 100 203 106
rect 145 23 149 100
rect 207 92 238 93
rect 159 89 238 92
rect 159 87 210 89
rect 159 81 164 87
rect 168 81 173 87
rect 205 81 210 87
rect 230 78 234 89
rect 305 78 313 169
rect 187 66 192 76
rect 228 73 313 78
rect 182 62 192 66
rect 236 66 241 73
rect 182 58 186 62
rect 248 66 253 73
rect 182 55 223 58
rect 182 52 186 55
rect 220 52 223 55
rect 263 52 268 61
rect 165 36 168 50
rect 210 47 212 50
rect 220 48 251 52
rect 263 48 417 52
rect 192 44 195 47
rect 209 36 212 47
rect 263 44 268 48
rect 165 31 212 36
rect 248 35 253 39
rect 269 35 277 36
rect 244 30 277 35
rect 269 29 277 30
rect 145 22 175 23
rect 145 19 180 22
rect 271 5 277 29
rect 10 0 277 5
rect -69 -30 443 -25
rect -912 -133 -747 -127
rect -715 -150 -706 -64
rect -1089 -156 -706 -150
<< m2contact >>
rect 683 651 695 662
rect -1313 607 -1302 617
rect -927 605 -913 615
rect -1202 577 -1195 583
rect -1159 552 -1154 557
rect -1032 577 -1027 582
rect -1161 534 -1156 539
rect -1101 551 -1094 556
rect -1138 534 -1133 539
rect -1084 511 -1079 516
rect -1005 539 -998 546
rect -990 537 -985 544
rect -930 534 -925 539
rect -916 509 -911 514
rect -820 491 -803 502
rect -1164 383 -1159 388
rect -1205 354 -1198 360
rect -1162 330 -1157 335
rect -1035 355 -1030 360
rect -1164 312 -1159 317
rect -1102 326 -1096 332
rect -1141 312 -1136 317
rect -1009 317 -1000 322
rect -1087 289 -1082 294
rect -933 312 -928 317
rect -919 287 -914 292
rect -767 467 -755 478
rect -818 425 -807 440
rect -847 402 -836 413
rect 275 606 288 619
rect 603 607 610 615
rect 1230 638 1240 647
rect 798 622 806 629
rect 726 614 736 621
rect 744 602 754 610
rect 874 618 883 624
rect 1378 615 1388 625
rect 893 603 901 609
rect -649 486 -637 502
rect -609 423 -599 430
rect -573 421 -560 431
rect -672 406 -661 417
rect -430 404 -418 418
rect -286 412 -271 421
rect 499 535 504 540
rect 592 542 598 549
rect 546 525 553 532
rect 635 535 640 540
rect 730 543 736 550
rect 484 510 489 517
rect 507 510 512 517
rect 682 525 689 532
rect 781 537 786 542
rect 876 544 882 551
rect 828 527 835 534
rect 928 537 933 542
rect 1032 544 1039 552
rect 620 510 625 517
rect 643 510 648 517
rect 766 512 771 519
rect 789 512 794 519
rect 975 527 982 534
rect 1140 536 1145 541
rect 893 511 901 517
rect 913 512 918 519
rect 936 512 941 519
rect 1187 526 1194 533
rect 1276 536 1281 541
rect 1125 511 1130 518
rect 1148 511 1153 518
rect 1323 526 1330 533
rect 1422 538 1427 543
rect 1469 528 1476 535
rect 1569 538 1574 543
rect 1261 511 1266 518
rect 1284 511 1289 518
rect 1407 513 1412 520
rect 1430 513 1435 520
rect 1616 528 1623 535
rect 1554 513 1559 520
rect 1577 513 1582 520
rect 499 427 504 432
rect 605 435 610 441
rect 546 417 553 424
rect 643 427 648 432
rect 745 433 751 440
rect -815 375 -803 385
rect -737 376 -726 385
rect 444 397 450 404
rect 484 401 489 409
rect 507 402 512 409
rect -728 324 -721 330
rect -629 315 -624 320
rect -573 325 -567 330
rect -678 305 -671 312
rect -482 315 -477 320
rect -429 322 -422 328
rect -1244 192 -1236 198
rect -1227 170 -1220 176
rect -1032 170 -1027 175
rect -1160 143 -1155 149
rect -1161 127 -1156 132
rect -1241 111 -1235 117
rect -1202 111 -1196 116
rect -1162 99 -1157 105
rect -1245 87 -1237 93
rect -1100 142 -1095 147
rect -1138 127 -1133 132
rect -1084 104 -1079 109
rect -1005 132 -997 137
rect -930 127 -925 132
rect -916 102 -911 107
rect -846 276 -834 287
rect -816 282 -805 292
rect -637 290 -632 297
rect -614 290 -609 297
rect -531 305 -524 312
rect -336 313 -331 318
rect -285 320 -279 325
rect -490 290 -485 297
rect -385 303 -378 310
rect -200 313 -195 318
rect -467 290 -462 297
rect -344 288 -339 295
rect -321 288 -316 295
rect -249 303 -242 310
rect -208 288 -203 295
rect -185 288 -180 295
rect -847 220 -837 233
rect -853 193 -843 201
rect -753 217 -747 222
rect -768 168 -758 178
rect -887 69 -878 76
rect -886 40 -879 47
rect -1202 -5 -1195 1
rect -1032 -5 -1027 0
rect -1160 -31 -1155 -26
rect -1161 -48 -1156 -43
rect -1100 -33 -1094 -28
rect -1138 -48 -1133 -43
rect -1010 -43 -1000 -38
rect -1084 -71 -1079 -66
rect -930 -48 -925 -43
rect -916 -73 -911 -68
rect -771 -61 -762 -49
rect -912 -118 -903 -108
rect 192 357 197 362
rect 272 366 278 371
rect 690 417 697 424
rect 792 429 797 434
rect 894 436 900 442
rect 839 419 846 426
rect 937 430 942 435
rect 1019 436 1027 443
rect 984 420 991 427
rect 628 402 633 409
rect 651 402 656 409
rect 777 404 782 411
rect 800 404 805 411
rect 922 404 927 411
rect 945 405 950 412
rect 239 348 246 354
rect 100 326 108 334
rect 177 333 182 340
rect 268 345 277 354
rect 444 362 450 367
rect 200 334 205 340
rect -726 215 -720 221
rect -638 208 -633 213
rect -584 217 -579 222
rect -687 198 -680 205
rect -493 207 -488 212
rect -443 213 -436 218
rect -646 183 -641 190
rect -623 182 -618 189
rect -542 197 -535 204
rect -344 205 -339 210
rect -298 214 -293 219
rect 17 227 22 232
rect 41 227 47 232
rect 54 227 59 232
rect 77 227 85 232
rect -501 182 -496 189
rect -478 182 -473 189
rect -393 195 -386 202
rect -200 205 -195 210
rect -352 180 -347 187
rect -329 180 -324 187
rect -249 195 -242 202
rect -208 180 -203 187
rect -185 179 -180 187
rect -144 179 -139 185
rect -70 179 -65 185
rect 53 205 59 210
rect -69 15 -62 21
rect 332 347 341 356
rect 191 239 196 244
rect 236 230 244 235
rect 176 214 181 219
rect 198 213 204 219
rect 282 144 290 150
rect 190 135 195 140
rect 235 126 243 132
rect 190 39 195 44
rect 417 47 427 54
rect 236 29 244 35
rect 198 15 203 22
rect 443 -33 451 -20
rect -717 -64 -703 -49
rect -1100 -156 -1089 -145
<< metal2 >>
rect 537 687 544 688
rect 537 686 805 687
rect 537 682 806 686
rect 537 653 544 682
rect 224 647 544 653
rect 567 661 572 662
rect 567 655 683 661
rect -1210 613 -1154 614
rect -1302 608 -1154 613
rect -1302 607 -1204 608
rect -1202 360 -1199 577
rect -1159 557 -1154 608
rect -1024 605 -927 611
rect -1024 602 -917 605
rect -1024 582 -1019 602
rect -1027 577 -1005 582
rect -1156 534 -1138 539
rect -1100 434 -1095 551
rect -1011 539 -1005 577
rect -998 539 -990 544
rect -930 539 -925 602
rect -1084 469 -1079 511
rect -926 509 -916 513
rect -926 469 -920 509
rect 225 506 233 647
rect 567 633 572 655
rect 800 660 806 682
rect -803 491 -649 499
rect -586 496 233 506
rect -1084 468 -778 469
rect -1084 464 -776 468
rect -755 473 -668 474
rect -755 467 -667 473
rect -931 463 -776 464
rect -792 461 -776 463
rect -1100 429 -818 434
rect -1202 203 -1199 354
rect -1162 335 -1159 383
rect -1027 380 -920 389
rect -1027 360 -1022 380
rect -1030 355 -1008 360
rect -1159 312 -1141 317
rect -1101 227 -1097 326
rect -1014 322 -1008 355
rect -1014 317 -1009 322
rect -933 317 -928 380
rect -1087 247 -1082 289
rect -929 287 -919 291
rect -846 287 -840 402
rect -813 292 -808 375
rect -929 247 -923 287
rect -1087 244 -923 247
rect -1087 242 -823 244
rect -934 241 -823 242
rect -1101 223 -847 227
rect -1227 199 -1199 203
rect -1227 198 -1224 199
rect -1236 192 -1224 198
rect -1160 196 -1156 197
rect -1227 176 -1224 192
rect -1188 193 -1156 196
rect -1188 181 -1183 193
rect -1202 178 -1183 181
rect -1242 111 -1241 116
rect -1242 93 -1239 111
rect -1227 93 -1224 170
rect -1202 116 -1198 178
rect -1160 149 -1156 193
rect -1024 195 -917 204
rect -1024 175 -1019 195
rect -1027 170 -1005 175
rect -1156 127 -1138 132
rect -1227 89 -1199 93
rect -1202 1 -1199 89
rect -1160 -26 -1157 99
rect -1099 44 -1095 142
rect -1011 132 -1005 170
rect -930 132 -925 195
rect -1084 62 -1079 104
rect -926 102 -916 106
rect -926 62 -920 102
rect -851 74 -846 193
rect -828 172 -823 241
rect -878 71 -846 74
rect -878 70 -847 71
rect -1084 60 -920 62
rect -830 61 -823 172
rect -788 134 -778 461
rect -672 417 -667 467
rect -607 407 -601 423
rect -608 383 -601 407
rect -726 376 -601 383
rect -768 331 -732 332
rect -768 330 -724 331
rect -768 326 -728 330
rect -768 178 -760 326
rect -755 325 -728 326
rect -655 315 -629 318
rect -655 311 -650 315
rect -671 306 -650 311
rect -585 295 -578 496
rect 225 495 233 496
rect 247 625 572 633
rect 591 629 768 634
rect 800 629 805 660
rect 1240 638 1241 647
rect 858 629 1068 634
rect 591 628 618 629
rect 247 485 253 625
rect -445 478 254 485
rect -573 330 -569 421
rect -508 315 -482 318
rect -508 311 -503 315
rect -524 306 -503 311
rect -609 292 -578 295
rect -609 291 -581 292
rect -637 272 -632 290
rect -490 272 -485 290
rect -445 294 -438 478
rect 276 456 282 606
rect 592 549 598 628
rect 730 621 735 622
rect 504 535 530 538
rect 525 531 530 535
rect 525 526 546 531
rect -296 448 282 456
rect 384 505 389 507
rect 484 506 489 510
rect 467 505 489 506
rect 384 501 489 505
rect 384 500 473 501
rect -429 328 -425 404
rect -362 313 -336 316
rect -362 309 -357 313
rect -378 304 -357 309
rect -462 290 -438 294
rect -467 289 -440 290
rect -296 291 -291 448
rect -135 434 -128 435
rect 384 434 389 500
rect 507 494 512 510
rect 603 514 608 607
rect 730 550 735 614
rect 763 602 768 629
rect 858 602 862 629
rect 640 535 666 538
rect 661 531 666 535
rect 661 526 682 531
rect 603 510 620 514
rect 746 515 751 602
rect 763 598 862 602
rect 876 551 881 618
rect 786 537 812 540
rect 807 533 812 537
rect 807 528 828 533
rect 746 512 766 515
rect 746 511 771 512
rect 751 510 767 511
rect 603 509 617 510
rect 603 508 608 509
rect 643 494 648 510
rect 789 494 794 512
rect 893 517 897 603
rect 1033 552 1039 599
rect 933 537 959 540
rect 954 533 959 537
rect 954 528 975 533
rect 901 515 909 516
rect 901 512 913 515
rect 901 511 918 512
rect 936 494 941 512
rect 1062 506 1068 629
rect 1145 536 1171 539
rect 1166 532 1171 536
rect 1166 527 1187 532
rect 1125 506 1130 511
rect 1062 501 1130 506
rect 1237 515 1241 638
rect 1388 615 1389 624
rect 1281 536 1307 539
rect 1302 532 1307 536
rect 1302 527 1323 532
rect 1236 511 1261 515
rect 1383 517 1389 615
rect 1527 597 1528 604
rect 1427 538 1453 541
rect 1448 534 1453 538
rect 1448 529 1469 534
rect 1383 516 1401 517
rect 1383 513 1407 516
rect 1383 512 1412 513
rect 1523 516 1528 597
rect 1574 538 1600 541
rect 1595 534 1600 538
rect 1595 529 1616 534
rect -135 428 389 434
rect -285 325 -279 412
rect -226 313 -200 316
rect -226 309 -221 313
rect -242 304 -221 309
rect -316 288 -290 291
rect -344 272 -339 288
rect -208 272 -203 288
rect -135 290 -128 428
rect 384 426 389 428
rect 422 491 941 494
rect 422 380 426 491
rect 504 427 530 430
rect 525 423 530 427
rect 605 424 610 435
rect 1027 438 1068 443
rect 648 427 674 430
rect 525 418 546 423
rect 669 423 674 427
rect 669 418 690 423
rect 745 412 751 433
rect 797 429 823 432
rect 818 425 823 429
rect 818 420 839 425
rect 896 414 900 436
rect 942 430 968 433
rect 963 426 968 430
rect 963 421 984 426
rect 473 404 484 405
rect 450 401 484 404
rect 507 380 512 402
rect 622 402 628 405
rect 622 401 633 402
rect 651 380 656 402
rect 771 404 777 407
rect 771 403 782 404
rect 800 380 805 404
rect 918 404 922 408
rect 945 380 950 405
rect 422 377 950 380
rect 278 367 295 371
rect 422 370 426 377
rect 945 376 950 377
rect 418 367 426 370
rect 197 357 223 360
rect 218 353 223 357
rect 218 349 239 353
rect 218 348 230 349
rect -180 288 -128 290
rect -185 285 -128 288
rect 45 326 100 331
rect 177 331 182 333
rect 108 326 182 331
rect -637 269 -118 272
rect -747 217 -726 221
rect -664 208 -638 211
rect -584 212 -581 217
rect -664 204 -659 208
rect -519 207 -493 210
rect -680 199 -659 204
rect -519 203 -514 207
rect -535 198 -514 203
rect -443 205 -440 213
rect -370 205 -344 208
rect -370 201 -365 205
rect -386 196 -365 201
rect -298 194 -294 214
rect -226 205 -200 208
rect -226 201 -221 205
rect -242 196 -221 201
rect -646 158 -641 183
rect -618 183 -596 187
rect -501 158 -496 182
rect -473 182 -457 184
rect -478 180 -457 182
rect -324 180 -314 184
rect -352 158 -347 180
rect -208 158 -203 180
rect -180 179 -144 183
rect -122 158 -118 269
rect 45 234 50 326
rect 200 316 205 334
rect 132 309 205 316
rect 45 232 49 234
rect 132 232 139 309
rect 196 239 219 242
rect 0 227 17 232
rect 47 227 49 232
rect 85 227 139 232
rect 214 235 219 239
rect 223 235 228 348
rect 277 348 332 354
rect 214 230 236 235
rect 0 201 6 227
rect 54 210 58 227
rect 132 215 139 227
rect 132 214 176 215
rect 132 208 181 214
rect 198 201 204 213
rect 0 197 204 201
rect 0 196 6 197
rect -646 155 -118 158
rect -646 154 -641 155
rect -788 131 -298 134
rect -788 130 -778 131
rect -492 110 -488 115
rect -493 107 -442 110
rect -435 107 -434 110
rect -493 106 -434 107
rect -616 92 -583 95
rect -616 91 -578 92
rect -830 60 -772 61
rect -492 60 -488 106
rect -308 76 -141 82
rect -1084 57 -837 60
rect -1099 40 -886 44
rect -1024 20 -917 29
rect -1024 0 -1019 20
rect -1027 -5 -1005 0
rect -1156 -48 -1138 -43
rect -1100 -128 -1096 -33
rect -1011 -38 -1005 -5
rect -1011 -43 -1010 -38
rect -930 -43 -925 20
rect -1084 -113 -1079 -71
rect -926 -73 -916 -69
rect -926 -112 -920 -73
rect -927 -113 -912 -112
rect -1084 -118 -912 -113
rect -846 -114 -837 57
rect -830 57 -485 60
rect -830 54 -772 57
rect -448 60 -170 62
rect -448 56 -169 60
rect -588 28 -206 32
rect -762 -61 -717 -52
rect -639 -112 -629 -111
rect -757 -113 -629 -112
rect -817 -114 -629 -113
rect -846 -117 -629 -114
rect -846 -118 -639 -117
rect -211 -108 -206 28
rect -179 -75 -169 56
rect -146 55 -141 76
rect -146 -23 -140 55
rect -122 -6 -118 155
rect -69 21 -66 179
rect 40 15 44 197
rect 195 135 219 138
rect 214 131 219 135
rect 223 131 228 230
rect 281 144 282 148
rect 290 144 331 148
rect 214 126 235 131
rect 195 39 218 42
rect 214 35 218 39
rect 223 35 228 126
rect 214 30 236 35
rect 40 12 203 15
rect 198 11 203 12
rect 325 -6 331 144
rect 418 54 422 367
rect 766 366 770 367
rect 446 339 449 362
rect -122 -11 331 -6
rect 325 -12 331 -11
rect 445 -20 449 339
rect 618 302 622 337
rect 766 312 770 360
rect 976 315 979 370
rect 1148 334 1153 511
rect 1284 349 1289 511
rect 1430 365 1435 513
rect 1522 513 1554 516
rect 1522 512 1559 513
rect 1577 495 1582 513
rect 1578 446 1582 495
rect 504 293 622 302
rect 765 303 770 312
rect 789 310 979 315
rect -145 -51 -140 -23
rect 504 -51 509 293
rect 531 263 540 265
rect 765 263 769 303
rect 531 255 772 263
rect -145 -57 514 -51
rect -179 -80 -170 -75
rect 531 -80 540 255
rect 789 241 801 310
rect 578 229 801 241
rect -179 -90 542 -80
rect 531 -92 540 -90
rect 579 -108 589 229
rect -211 -117 589 -108
rect -1100 -145 -1095 -128
<< m3contact >>
rect 1033 599 1041 607
rect 1518 597 1527 607
rect 1068 436 1078 444
rect 605 418 610 424
rect 616 399 622 407
rect 744 405 751 412
rect 765 400 771 408
rect 895 407 901 414
rect 910 402 918 412
rect 973 370 980 376
rect -584 207 -579 212
rect -443 200 -438 205
rect -298 189 -293 194
rect -596 183 -591 189
rect -457 179 -450 185
rect -314 180 -308 187
rect -298 130 -293 135
rect -442 107 -435 113
rect -625 90 -616 98
rect -583 92 -576 98
rect -316 76 -308 86
rect -457 56 -448 65
rect -593 28 -588 36
rect -629 -120 -617 -107
rect 765 360 772 366
rect 616 337 624 344
rect 1577 437 1587 446
rect 1428 357 1438 365
rect 1281 342 1291 349
rect 1148 326 1155 334
<< metal3 >>
rect 1041 605 1051 606
rect 1041 600 1518 605
rect 1041 599 1051 600
rect 1073 444 1577 446
rect 1078 437 1577 444
rect 605 329 610 418
rect 617 344 622 399
rect 744 349 751 405
rect 766 366 770 400
rect 895 362 901 407
rect 912 374 915 402
rect 912 371 973 374
rect 895 357 1428 362
rect 744 343 1281 349
rect 605 326 1148 329
rect 605 325 1154 326
rect -591 183 -590 188
rect -627 90 -625 96
rect -627 -107 -622 90
rect -593 36 -590 183
rect -582 98 -579 207
rect -457 65 -451 179
rect -442 113 -439 200
rect -315 180 -314 182
rect -315 86 -309 180
rect -298 135 -294 189
<< labels >>
rlabel metal1 38 230 38 230 1 S0c
rlabel metal1 23 230 23 230 1 S0
rlabel metal1 61 231 61 231 1 S1
rlabel metal1 277 250 277 250 1 D1
rlabel metal1 271 369 271 369 1 D0
rlabel metal1 279 50 279 50 1 D3
rlabel metal1 188 33 188 33 1 DEC_AND_NODE_4
rlabel metal1 188 56 188 56 1 DEC_D3_NAND
rlabel metal1 280 146 280 146 1 D2
rlabel metal1 189 129 189 129 1 DEC_AND_NODE_3
rlabel metal1 189 152 189 152 1 DEC_D2_NAND
rlabel metal1 191 233 191 233 1 Dec_AND_node_2
rlabel metal1 192 256 192 256 1 DEC_D1_NAND
rlabel metal1 187 375 187 375 1 DEC_D0_NAND
rlabel metal1 192 352 192 352 1 Dec_AND_node_1
rlabel m2contact 80 230 80 230 1 S1c
rlabel metal1 80 212 80 212 1 gnd
rlabel metal1 56 256 56 256 1 vdd
rlabel metal2 479 403 479 403 1 B3
rlabel m3contact 620 404 620 404 1 B2
rlabel metal2 772 406 772 406 1 B1
rlabel metal1 938 424 938 424 1 ander_node_5
rlabel metal1 790 424 790 424 1 ander_node_6
rlabel metal1 641 420 641 420 1 ander_node_7
rlabel metal1 496 422 496 422 1 ander_node_8
rlabel metal1 972 441 972 441 1 and_b0e_nand
rlabel metal1 837 440 837 440 1 and_b1e_nand
rlabel metal1 683 437 683 437 1 and_b2e_nand
rlabel metal1 535 437 535 437 1 and_b3e_nand
rlabel metal1 1016 441 1016 441 1 and_b0e
rlabel metal1 872 440 872 440 1 and_b1e
rlabel metal1 724 437 724 437 1 and_b2e
rlabel metal1 580 438 580 438 1 and_b3e
rlabel metal1 1007 547 1007 547 1 and_a0e
rlabel metal1 860 547 860 547 1 and_a1e
rlabel metal1 713 545 713 545 1 and_a2e
rlabel metal1 578 546 578 546 1 and_a3e
rlabel metal1 970 547 970 547 1 and_a0e_nand
rlabel metal1 824 548 824 548 1 and_a1e_nand
rlabel metal1 681 546 681 546 1 and_a2e_nand
rlabel metal1 537 547 537 547 1 and_a3e_nand
rlabel metal1 927 531 927 531 1 ander_node_4
rlabel metal1 780 531 780 531 1 ander_node_3
rlabel metal1 634 530 634 530 1 ander_node_2
rlabel metal1 498 529 498 529 1 ander_node_1
rlabel metal2 907 513 907 513 1 A0
rlabel metal2 761 513 761 513 1 A1
rlabel metal2 614 511 614 511 1 A2
rlabel metal2 486 506 486 506 1 A3
rlabel metal1 1138 531 1138 531 1 ander_node_9
rlabel metal1 1272 531 1272 531 1 ander_node_10
rlabel metal1 1422 534 1422 534 1 ander_node_11
rlabel metal1 1566 531 1566 531 1 ander_node_12
rlabel metal1 1179 547 1179 547 1 A3_and_B3_nand
rlabel metal1 1307 548 1307 548 1 A2_and_B2_nand
rlabel metal1 1462 549 1462 549 1 A1_and_B1_nand
rlabel metal1 1602 549 1602 549 1 A0_and_B0_nand
rlabel metal1 1220 547 1220 547 1 A3_and_B3
rlabel metal1 1356 547 1356 547 1 A2_and_B2
rlabel metal1 1501 549 1501 549 1 A1_and_B1
rlabel metal1 1649 549 1649 549 1 A0_and_B0
rlabel metal1 -191 308 -191 308 1 compare_node_1
rlabel metal1 -330 308 -330 308 1 compare_node_2
rlabel metal1 -476 309 -476 309 1 compare_node_3
rlabel metal1 -622 309 -622 309 1 compare_node_4
rlabel metal1 -631 203 -631 203 1 compare_node_5
rlabel metal1 -487 201 -487 201 1 compare_node_6
rlabel metal1 -337 198 -337 198 1 compare_node_7
rlabel metal1 -194 198 -194 198 1 compare_node_8
rlabel metal1 -191 339 -191 339 1 compare_A3e_nand
rlabel metal1 -325 338 -325 338 1 compare_A2e_nand
rlabel metal1 -471 337 -471 337 1 compare_A1e_nand
rlabel metal1 -619 341 -619 341 1 compare_A0e_nand
rlabel metal1 -627 234 -627 234 1 compare_B0e_nand
rlabel metal1 -482 231 -482 231 1 compare_B1e_nand
rlabel metal1 -334 230 -334 230 1 compare_B2e_nand
rlabel metal1 -189 230 -189 230 1 compare_B3e_nand
rlabel metal1 -275 324 -275 324 1 compare_A3e
rlabel metal1 -410 325 -410 325 1 compare_A2e
rlabel metal1 -554 325 -554 325 1 compare_A1e
rlabel metal1 -703 327 -703 327 1 compare_A0e
rlabel metal1 -711 219 -711 219 1 compare_B0e
rlabel metal1 -565 218 -565 218 1 compare_B1e
rlabel metal1 -416 215 -416 215 1 compare_B2e
rlabel metal1 -271 216 -271 216 1 compare_B3e
rlabel pdiffusion -1053 564 -1053 564 1 xnor_1
rlabel ndiffusion -1053 524 -1053 524 1 xnor_2
rlabel metal1 -992 553 -992 553 1 xor_1
rlabel ndiffusion -971 564 -971 564 1 xnor_3
rlabel pdiffusion -971 524 -971 524 1 xnor_4
rlabel metal1 -963 478 -963 478 1 A3c
rlabel metal1 -1006 595 -1006 595 1 B3c
rlabel pdiffusion -1058 342 -1058 342 1 xnor_5
rlabel ndiffusion -1055 302 -1055 302 1 xnor_6
rlabel ndiffusion -972 342 -972 342 1 xnor_7
rlabel pdiffusion -976 301 -976 301 1 xnor_8
rlabel metal1 -964 253 -964 253 1 A2c
rlabel metal1 -1005 375 -1005 375 1 B2c
rlabel metal1 -1005 190 -1005 190 1 B1c
rlabel metal1 -971 67 -971 67 1 A1c
rlabel pdiffusion -1053 156 -1053 156 1 xnor_9
rlabel ndiffusion -1050 117 -1050 117 1 xnor_10
rlabel pdiffusion -972 117 -972 117 1 xnor_11
rlabel ndiffusion -970 157 -970 157 1 xnor_12
rlabel metal1 -1003 329 -1003 329 1 xor_2
rlabel metal1 -998 145 -998 145 1 xor_3
rlabel metal1 -995 14 -995 14 1 B0c
rlabel metal1 -971 -107 -971 -107 1 A0c
rlabel metal1 -995 -29 -995 -29 1 xor_4
rlabel pdiffusion -1054 -18 -1054 -18 1 xnor_13
rlabel ndiffusion -1052 -59 -1052 -59 1 xnor_14
rlabel ndiffusion -970 -19 -970 -19 1 xnor_15
rlabel pdiffusion -970 -58 -970 -58 1 xnor_16
rlabel ndiffusion -1300 134 -1300 134 1 A_compare_B_node_3
rlabel ndiffusion -1283 135 -1283 135 1 A_compare_B_node_2
rlabel ndiffusion -1268 135 -1268 135 1 A_compare_B_node_1
rlabel metal1 -1383 159 -1383 159 3 A_equal_B
rlabel metal1 -1337 147 -1337 147 1 A_equal_B_c
rlabel metal1 -1294 217 -1294 217 1 A2e_xnor_B2e
rlabel metal1 -1165 555 -1165 555 1 A3e_xnor_B3e
rlabel metal1 -1166 147 -1166 147 1 A1e_xnor_B1e
rlabel metal1 -1165 -29 -1165 -29 1 A0e_xnor_B0e
rlabel metal2 919 405 919 405 1 B0
<< end >>
