magic
tech scmos
timestamp 1699124852
<< nwell >>
rect -35 -6 42 26
<< ntransistor >>
rect -20 -25 -15 -20
rect -4 -25 1 -20
rect 12 -25 17 -20
<< ptransistor >>
rect -20 9 -15 14
rect -4 9 1 14
rect 12 9 17 14
<< ndiffusion >>
rect -23 -25 -20 -20
rect -15 -25 -4 -20
rect 1 -25 12 -20
rect 17 -25 23 -20
<< pdiffusion >>
rect -23 9 -20 14
rect -15 9 -12 14
rect -7 9 -4 14
rect 1 9 4 14
rect 9 9 12 14
rect 17 9 20 14
<< ndcontact >>
rect -28 -25 -23 -20
rect 23 -25 28 -20
<< pdcontact >>
rect -28 9 -23 14
rect -12 9 -7 14
rect 4 9 9 14
rect 20 9 25 14
<< nsubstratencontact >>
rect 30 9 35 14
<< polysilicon >>
rect -20 14 -15 19
rect -4 14 1 19
rect 12 14 17 19
rect -20 -9 -15 9
rect -4 -9 1 9
rect 12 -9 17 9
rect -19 -14 -15 -9
rect -3 -14 1 -9
rect 13 -14 17 -9
rect -20 -20 -15 -14
rect -4 -20 1 -14
rect 12 -20 17 -14
rect -20 -29 -15 -25
rect -4 -29 1 -25
rect 12 -29 17 -25
<< polycontact >>
rect -24 -14 -19 -9
rect -8 -14 -3 -9
rect 8 -14 13 -9
<< metal1 >>
rect -35 26 42 31
rect -28 14 -23 26
rect 4 14 9 26
rect 30 14 35 26
rect 25 9 26 14
rect -12 6 -7 9
rect 20 6 26 9
rect -12 1 26 6
rect 45 1 60 5
rect 83 1 88 5
rect -26 -14 -24 -9
rect -10 -14 -8 -9
rect 6 -14 8 -9
rect 23 -12 28 1
rect 45 -12 49 1
rect 23 -17 49 -12
rect 23 -20 28 -17
rect -28 -32 -23 -25
rect 52 -32 57 -12
rect -28 -36 57 -32
use not_without_labels  not_without_labels_0
timestamp 1699100137
transform 1 0 58 0 1 -5
box -16 -12 33 36
<< labels >>
rlabel metal1 -25 -11 -25 -11 1 input_A
rlabel metal1 -9 -11 -9 -11 1 input_B
rlabel metal1 7 -12 7 -12 1 input_C
rlabel ndiffusion 8 -22 8 -22 1 node_1
rlabel ndiffusion -9 -22 -9 -22 1 node_2
rlabel metal1 21 4 21 4 1 v_output_nand_3
rlabel metal1 -2 28 -2 28 5 Vdd!
rlabel metal1 -25 -26 -25 -26 1 Gnd!
rlabel metal1 87 2 87 2 7 v_output_and_3
<< end >>
