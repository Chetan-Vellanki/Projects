magic
tech scmos
timestamp 1701343358
<< nwell >>
rect 0 50 61 67
rect 75 34 121 53
rect 136 50 197 67
rect 211 34 257 53
rect 282 52 343 69
rect 357 36 403 55
rect 429 52 490 69
rect 504 36 550 55
rect 0 -58 61 -41
rect 75 -74 121 -55
rect 144 -58 205 -41
rect 219 -74 265 -55
rect 293 -56 354 -39
rect 368 -72 414 -53
rect 438 -55 499 -38
rect 513 -71 559 -52
<< ntransistor >>
rect 20 27 25 32
rect 43 27 48 32
rect 156 27 161 32
rect 179 27 184 32
rect 302 29 307 34
rect 325 29 330 34
rect 101 19 106 24
rect 237 19 242 24
rect 449 29 454 34
rect 472 29 477 34
rect 383 21 388 26
rect 530 21 535 26
rect 20 -81 25 -76
rect 43 -81 48 -76
rect 164 -81 169 -76
rect 187 -81 192 -76
rect 313 -79 318 -74
rect 336 -79 341 -74
rect 458 -78 463 -73
rect 481 -78 486 -73
rect 101 -89 106 -84
rect 245 -89 250 -84
rect 394 -87 399 -82
rect 539 -86 544 -81
<< ptransistor >>
rect 20 56 25 61
rect 43 56 48 61
rect 156 56 161 61
rect 179 56 184 61
rect 302 58 307 63
rect 325 58 330 63
rect 449 58 454 63
rect 472 58 477 63
rect 101 41 106 46
rect 237 41 242 46
rect 383 43 388 48
rect 530 43 535 48
rect 20 -52 25 -47
rect 43 -52 48 -47
rect 164 -52 169 -47
rect 187 -52 192 -47
rect 313 -50 318 -45
rect 336 -50 341 -45
rect 458 -49 463 -44
rect 481 -49 486 -44
rect 101 -67 106 -62
rect 245 -67 250 -62
rect 394 -65 399 -60
rect 539 -64 544 -59
<< ndiffusion >>
rect 18 27 20 32
rect 25 27 27 32
rect 41 27 43 32
rect 48 27 50 32
rect 154 27 156 32
rect 161 27 163 32
rect 177 27 179 32
rect 184 27 186 32
rect 300 29 302 34
rect 307 29 309 34
rect 323 29 325 34
rect 330 29 332 34
rect 99 19 101 24
rect 106 19 109 24
rect 235 19 237 24
rect 242 19 245 24
rect 447 29 449 34
rect 454 29 456 34
rect 470 29 472 34
rect 477 29 479 34
rect 381 21 383 26
rect 388 21 391 26
rect 528 21 530 26
rect 535 21 538 26
rect 18 -81 20 -76
rect 25 -81 27 -76
rect 41 -81 43 -76
rect 48 -81 50 -76
rect 162 -81 164 -76
rect 169 -81 171 -76
rect 185 -81 187 -76
rect 192 -81 194 -76
rect 311 -79 313 -74
rect 318 -79 320 -74
rect 334 -79 336 -74
rect 341 -79 343 -74
rect 456 -78 458 -73
rect 463 -78 465 -73
rect 479 -78 481 -73
rect 486 -78 488 -73
rect 99 -89 101 -84
rect 106 -89 109 -84
rect 243 -89 245 -84
rect 250 -89 253 -84
rect 392 -87 394 -82
rect 399 -87 402 -82
rect 537 -86 539 -81
rect 544 -86 547 -81
<< pdiffusion >>
rect 18 56 20 61
rect 25 56 32 61
rect 37 56 43 61
rect 48 56 50 61
rect 154 56 156 61
rect 161 56 168 61
rect 173 56 179 61
rect 184 56 186 61
rect 300 58 302 63
rect 307 58 314 63
rect 319 58 325 63
rect 330 58 332 63
rect 447 58 449 63
rect 454 58 461 63
rect 466 58 472 63
rect 477 58 479 63
rect 99 41 101 46
rect 106 41 109 46
rect 235 41 237 46
rect 242 41 245 46
rect 381 43 383 48
rect 388 43 391 48
rect 528 43 530 48
rect 535 43 538 48
rect 18 -52 20 -47
rect 25 -52 32 -47
rect 37 -52 43 -47
rect 48 -52 50 -47
rect 162 -52 164 -47
rect 169 -52 176 -47
rect 181 -52 187 -47
rect 192 -52 194 -47
rect 311 -50 313 -45
rect 318 -50 325 -45
rect 330 -50 336 -45
rect 341 -50 343 -45
rect 456 -49 458 -44
rect 463 -49 470 -44
rect 475 -49 481 -44
rect 486 -49 488 -44
rect 99 -67 101 -62
rect 106 -67 109 -62
rect 243 -67 245 -62
rect 250 -67 253 -62
rect 392 -65 394 -60
rect 399 -65 402 -60
rect 537 -64 539 -59
rect 544 -64 547 -59
<< ndcontact >>
rect 13 27 18 32
rect 27 27 31 32
rect 37 27 41 32
rect 50 27 55 32
rect 149 27 154 32
rect 163 27 167 32
rect 173 27 177 32
rect 186 27 191 32
rect 295 29 300 34
rect 309 29 313 34
rect 319 29 323 34
rect 332 29 337 34
rect 94 19 99 24
rect 109 19 114 24
rect 230 19 235 24
rect 245 19 250 24
rect 442 29 447 34
rect 456 29 460 34
rect 466 29 470 34
rect 479 29 484 34
rect 376 21 381 26
rect 391 21 396 26
rect 523 21 528 26
rect 538 21 543 26
rect 13 -81 18 -76
rect 27 -81 31 -76
rect 37 -81 41 -76
rect 50 -81 55 -76
rect 157 -81 162 -76
rect 171 -81 175 -76
rect 181 -81 185 -76
rect 194 -81 199 -76
rect 306 -79 311 -74
rect 320 -79 324 -74
rect 330 -79 334 -74
rect 343 -79 348 -74
rect 451 -78 456 -73
rect 465 -78 469 -73
rect 475 -78 479 -73
rect 488 -78 493 -73
rect 94 -89 99 -84
rect 109 -89 114 -84
rect 238 -89 243 -84
rect 253 -89 258 -84
rect 387 -87 392 -82
rect 402 -87 407 -82
rect 532 -86 537 -81
rect 547 -86 552 -81
<< pdcontact >>
rect 13 56 18 61
rect 32 56 37 61
rect 50 56 55 61
rect 149 56 154 61
rect 168 56 173 61
rect 186 56 191 61
rect 295 58 300 63
rect 314 58 319 63
rect 332 58 337 63
rect 442 58 447 63
rect 461 58 466 63
rect 479 58 484 63
rect 94 41 99 46
rect 109 41 114 46
rect 230 41 235 46
rect 245 41 250 46
rect 376 43 381 48
rect 391 43 396 48
rect 523 43 528 48
rect 538 43 543 48
rect 13 -52 18 -47
rect 32 -52 37 -47
rect 50 -52 55 -47
rect 157 -52 162 -47
rect 176 -52 181 -47
rect 194 -52 199 -47
rect 306 -50 311 -45
rect 325 -50 330 -45
rect 343 -50 348 -45
rect 451 -49 456 -44
rect 470 -49 475 -44
rect 488 -49 493 -44
rect 94 -67 99 -62
rect 109 -67 114 -62
rect 238 -67 243 -62
rect 253 -67 258 -62
rect 387 -65 392 -60
rect 402 -65 407 -60
rect 532 -64 537 -59
rect 547 -64 552 -59
<< nsubstratencontact >>
rect 4 56 9 61
rect 140 56 145 61
rect 286 58 291 63
rect 433 58 438 63
rect 82 41 87 46
rect 218 41 223 46
rect 364 43 369 48
rect 511 43 516 48
rect 4 -52 9 -47
rect 148 -52 153 -47
rect 297 -50 302 -45
rect 442 -49 447 -44
rect 82 -67 87 -62
rect 226 -67 231 -62
rect 375 -65 380 -60
rect 520 -64 525 -59
<< polysilicon >>
rect 20 61 25 75
rect 43 61 48 75
rect 156 61 161 75
rect 179 61 184 75
rect 302 63 307 77
rect 325 63 330 77
rect 449 63 454 77
rect 472 63 477 77
rect 20 32 25 56
rect 43 32 48 56
rect 101 46 106 49
rect 101 32 106 41
rect 156 32 161 56
rect 179 32 184 56
rect 237 46 242 49
rect 237 32 242 41
rect 302 34 307 58
rect 325 34 330 58
rect 383 48 388 51
rect 383 34 388 43
rect 449 34 454 58
rect 472 34 477 58
rect 530 48 535 51
rect 530 34 535 43
rect 102 28 106 32
rect 20 8 25 27
rect 43 8 48 27
rect 101 24 106 28
rect 238 28 242 32
rect 384 30 388 34
rect 101 14 106 19
rect 156 8 161 27
rect 179 8 184 27
rect 237 24 242 28
rect 237 14 242 19
rect 302 10 307 29
rect 325 10 330 29
rect 383 26 388 30
rect 531 30 535 34
rect 383 16 388 21
rect 449 10 454 29
rect 472 10 477 29
rect 530 26 535 30
rect 530 16 535 21
rect 20 -47 25 -33
rect 43 -47 48 -33
rect 164 -47 169 -33
rect 187 -47 192 -33
rect 313 -45 318 -31
rect 336 -45 341 -31
rect 458 -44 463 -30
rect 481 -44 486 -30
rect 20 -76 25 -52
rect 43 -76 48 -52
rect 101 -62 106 -59
rect 101 -76 106 -67
rect 164 -76 169 -52
rect 187 -76 192 -52
rect 245 -62 250 -59
rect 245 -76 250 -67
rect 313 -74 318 -50
rect 336 -74 341 -50
rect 394 -60 399 -57
rect 394 -74 399 -65
rect 458 -73 463 -49
rect 481 -73 486 -49
rect 539 -59 544 -56
rect 539 -73 544 -64
rect 102 -80 106 -76
rect 20 -100 25 -81
rect 43 -100 48 -81
rect 101 -84 106 -80
rect 246 -80 250 -76
rect 395 -78 399 -74
rect 540 -77 544 -73
rect 101 -94 106 -89
rect 164 -100 169 -81
rect 187 -100 192 -81
rect 245 -84 250 -80
rect 245 -94 250 -89
rect 313 -98 318 -79
rect 336 -98 341 -79
rect 394 -82 399 -78
rect 394 -92 399 -87
rect 458 -97 463 -78
rect 481 -97 486 -78
rect 539 -81 544 -77
rect 539 -91 544 -86
<< polycontact >>
rect 97 28 102 32
rect 20 2 25 8
rect 233 28 238 32
rect 379 30 384 34
rect 43 2 48 8
rect 156 2 161 8
rect 179 2 184 8
rect 302 4 307 10
rect 526 30 531 34
rect 325 4 330 10
rect 449 4 454 10
rect 472 4 477 10
rect 97 -80 102 -76
rect 20 -106 25 -100
rect 241 -80 246 -76
rect 390 -78 395 -74
rect 535 -77 540 -73
rect 43 -106 48 -100
rect 164 -106 169 -100
rect 187 -106 192 -100
rect 313 -104 318 -98
rect 336 -104 341 -98
rect 458 -103 463 -97
rect 481 -103 486 -97
<< metal1 >>
rect 334 74 434 75
rect 481 74 512 75
rect 286 73 512 74
rect 52 72 83 73
rect 188 72 512 73
rect -17 71 512 72
rect -17 69 337 71
rect -17 67 55 69
rect -17 66 10 67
rect -17 -34 -9 66
rect 4 61 9 66
rect 13 61 18 67
rect 50 61 55 67
rect 75 68 191 69
rect 75 58 79 68
rect 140 67 191 68
rect 140 61 145 67
rect 32 46 37 56
rect 75 53 123 58
rect 149 61 154 67
rect 186 61 191 67
rect 211 58 215 69
rect 286 63 291 69
rect 295 63 300 69
rect 332 63 337 69
rect 357 60 361 71
rect 433 69 484 71
rect 433 63 438 69
rect 27 42 37 46
rect 82 46 87 53
rect 27 38 31 42
rect 94 46 99 53
rect 168 46 173 56
rect 211 53 259 58
rect 27 35 68 38
rect 27 32 31 35
rect 65 32 68 35
rect 109 32 114 41
rect 163 42 173 46
rect 218 46 223 53
rect 163 38 167 42
rect 230 46 235 53
rect 314 48 319 58
rect 357 55 405 60
rect 442 63 447 69
rect 479 63 484 69
rect 504 60 508 71
rect 163 35 204 38
rect 163 32 167 35
rect 201 32 204 35
rect 245 32 250 41
rect 309 44 319 48
rect 364 48 369 55
rect 309 40 313 44
rect 376 48 381 55
rect 461 48 466 58
rect 504 55 552 60
rect 309 37 350 40
rect 309 34 313 37
rect 347 34 350 37
rect 391 34 396 43
rect 456 44 466 48
rect 511 48 516 55
rect 456 40 460 44
rect 523 48 528 55
rect 456 37 497 40
rect 456 34 460 37
rect 494 34 497 37
rect 538 34 543 43
rect 10 16 13 30
rect 55 27 57 30
rect 65 28 97 32
rect 109 28 117 32
rect 37 24 40 27
rect 54 16 57 27
rect 109 24 114 28
rect 10 11 57 16
rect 94 15 99 19
rect 146 16 149 30
rect 191 27 193 30
rect 201 28 233 32
rect 245 28 253 32
rect 173 24 176 27
rect 190 16 193 27
rect 245 24 250 28
rect 89 10 124 15
rect 146 11 193 16
rect 20 1 25 2
rect 43 1 48 2
rect 120 -11 124 10
rect 230 15 235 19
rect 292 18 295 32
rect 337 29 339 32
rect 347 30 379 34
rect 391 30 399 34
rect 319 26 322 29
rect 336 18 339 29
rect 391 26 396 30
rect 225 14 260 15
rect 225 10 273 14
rect 292 13 339 18
rect 376 17 381 21
rect 439 18 442 32
rect 484 29 486 32
rect 494 30 526 34
rect 538 30 546 34
rect 466 26 469 29
rect 483 18 486 29
rect 538 26 543 30
rect 371 12 409 17
rect 439 13 486 18
rect 254 9 273 10
rect 156 1 161 2
rect 179 1 184 2
rect 264 -11 271 9
rect 302 3 307 4
rect 325 3 330 4
rect 400 -11 409 12
rect 523 17 528 21
rect 518 12 554 17
rect 449 3 454 4
rect 472 3 477 4
rect 545 -11 554 12
rect 573 -11 581 -10
rect 120 -17 581 -11
rect 490 -33 521 -32
rect 345 -34 521 -33
rect -17 -36 13 -34
rect 221 -35 521 -34
rect 52 -36 83 -35
rect 196 -36 521 -35
rect -17 -37 493 -36
rect -17 -39 348 -37
rect 357 -38 493 -37
rect -17 -41 55 -39
rect 74 -41 199 -39
rect 4 -47 9 -41
rect 13 -47 18 -41
rect 50 -47 55 -41
rect 75 -50 79 -41
rect 148 -47 153 -41
rect 32 -62 37 -52
rect 75 -55 123 -50
rect 157 -47 162 -41
rect 194 -47 199 -41
rect 219 -50 223 -39
rect 297 -45 302 -39
rect 306 -45 311 -39
rect 343 -45 348 -39
rect 368 -48 372 -38
rect 442 -44 447 -38
rect 27 -66 37 -62
rect 82 -62 87 -55
rect 27 -70 31 -66
rect 94 -62 99 -55
rect 176 -62 181 -52
rect 219 -55 267 -50
rect 27 -73 68 -70
rect 27 -76 31 -73
rect 65 -76 68 -73
rect 109 -76 114 -67
rect 171 -66 181 -62
rect 226 -62 231 -55
rect 171 -70 175 -66
rect 238 -62 243 -55
rect 325 -60 330 -50
rect 368 -53 416 -48
rect 451 -44 456 -38
rect 488 -44 493 -38
rect 513 -47 517 -36
rect 171 -73 212 -70
rect 171 -76 175 -73
rect 209 -76 212 -73
rect 253 -76 258 -67
rect 320 -64 330 -60
rect 375 -60 380 -53
rect 320 -68 324 -64
rect 387 -60 392 -53
rect 470 -59 475 -49
rect 513 -52 561 -47
rect 320 -71 361 -68
rect 320 -74 324 -71
rect 358 -74 361 -71
rect 402 -74 407 -65
rect 465 -63 475 -59
rect 520 -59 525 -52
rect 465 -67 469 -63
rect 532 -59 537 -52
rect 465 -70 506 -67
rect 465 -73 469 -70
rect 503 -73 506 -70
rect 547 -73 552 -64
rect 10 -92 13 -78
rect 55 -81 57 -78
rect 65 -80 97 -76
rect 109 -80 117 -76
rect 37 -84 40 -81
rect 54 -92 57 -81
rect 109 -84 114 -80
rect 10 -97 57 -92
rect 94 -93 99 -89
rect 154 -92 157 -78
rect 199 -81 201 -78
rect 209 -80 241 -76
rect 253 -80 261 -76
rect 181 -84 184 -81
rect 198 -92 201 -81
rect 253 -84 258 -80
rect 89 -98 124 -93
rect 154 -97 201 -92
rect 20 -107 25 -106
rect 43 -107 48 -106
rect 116 -122 125 -98
rect 238 -93 243 -89
rect 303 -90 306 -76
rect 348 -79 350 -76
rect 358 -78 390 -74
rect 402 -78 410 -74
rect 330 -82 333 -79
rect 347 -90 350 -79
rect 402 -82 407 -78
rect 233 -98 274 -93
rect 303 -95 350 -90
rect 387 -91 392 -87
rect 448 -89 451 -75
rect 493 -78 495 -75
rect 503 -77 535 -73
rect 547 -77 555 -73
rect 475 -81 478 -78
rect 492 -89 495 -78
rect 547 -81 552 -77
rect 382 -96 417 -91
rect 448 -94 495 -89
rect 532 -90 537 -86
rect 556 -90 563 -89
rect 527 -95 563 -90
rect 164 -107 169 -106
rect 187 -107 192 -106
rect 266 -122 273 -98
rect 313 -105 318 -104
rect 336 -105 341 -104
rect 410 -122 417 -96
rect 458 -105 463 -103
rect 481 -104 486 -103
rect 556 -122 563 -95
rect 116 -123 563 -122
rect 573 -123 581 -17
rect 116 -128 581 -123
rect 266 -130 273 -128
rect 556 -129 563 -128
<< m2contact >>
rect 35 19 40 24
rect 82 9 89 16
rect 171 19 176 24
rect 20 -6 25 1
rect 43 -6 48 1
rect 218 9 225 16
rect 317 21 322 26
rect 364 11 371 18
rect 464 21 469 26
rect 156 -6 161 1
rect 179 -6 184 1
rect 302 -4 307 3
rect 325 -4 330 3
rect 511 11 518 18
rect 449 -4 454 3
rect 472 -4 477 3
rect 35 -89 40 -84
rect 82 -99 89 -92
rect 179 -89 184 -84
rect 20 -115 25 -107
rect 43 -114 48 -107
rect 226 -99 233 -92
rect 328 -87 333 -82
rect 375 -97 382 -90
rect 473 -86 478 -81
rect 520 -96 527 -89
rect 164 -114 169 -107
rect 187 -114 192 -107
rect 313 -112 318 -105
rect 336 -112 341 -105
rect 458 -112 463 -105
rect 481 -111 486 -104
<< metal2 >>
rect 40 19 66 22
rect 176 19 202 22
rect 322 21 348 24
rect 469 21 495 24
rect 61 15 66 19
rect 61 10 82 15
rect 197 15 202 19
rect 343 17 348 21
rect 197 10 218 15
rect 343 12 364 17
rect 490 17 495 21
rect 490 12 511 17
rect 43 -22 48 -6
rect 179 -22 184 -6
rect 325 -22 330 -4
rect 472 -22 477 -4
rect -42 -25 477 -22
rect -42 -136 -38 -25
rect 40 -89 66 -86
rect 184 -89 210 -86
rect 333 -87 359 -84
rect 478 -86 504 -83
rect 61 -93 66 -89
rect 61 -98 82 -93
rect 205 -93 210 -89
rect 354 -91 359 -87
rect 499 -90 504 -86
rect 205 -98 226 -93
rect 354 -96 375 -91
rect 499 -95 520 -90
rect 43 -136 48 -114
rect 187 -136 192 -114
rect 336 -136 341 -112
rect 481 -136 486 -111
rect -42 -139 486 -136
rect 481 -140 486 -139
<< end >>
