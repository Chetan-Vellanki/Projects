* SPICE3 file created from DEC_AND_COMPARE.ext - technology: scmos

.option scale=90n

M1000 A_greater_B_node_8 A3e_xnor_B3e A_greater_B_node_9 Gnd nfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1001 and_b1e_nand B1 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1002 Dec_AND_node_1 S1c gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1003 and_a1e_nand A1 ander_node_3 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1004 xor_2 B2c xnor_7 Gnd nfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1005 vdd D3 and_b1e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1006 vdd A1 compare_A1e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1007 B0c compare_B0e gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1008 gnd A_equal_B_c A_LS_B_node_1 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1009 xor_1 B3c xnor_1 vdd pfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1010 ander_node_3 D3 gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1011 xor_4 A0c xnor_16 vdd pfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1012 A_greater_B_node_3 compare_A2e A3_eq_B3_A2_gt_B2_c Gnd nfet w=5 l=5
+  ad=27p pd=16u as=55p ps=32u
M1013 B3c compare_B3e vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1014 gnd compare_B3e_nand compare_B3e Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1015 gnd A3_eq_B3_A2_gt_B2_c A3_eq_B3_A2_gt_B2 Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1016 vdd D3 and_a2e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1017 A0_and_B0 A0_and_B0_nand vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1018 and_b2e_nand B2 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1019 B2c compare_B2e vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1020 and_a3e_nand A3 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1021 and_a3e and_a3e_nand vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1022 A_compare_B_node_2 A2e_xnor_B2e A_compare_B_node_3 Gnd nfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1023 and_a2e_nand A2 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1024 vdd A0e_xnor_B0e A_equal_B_c vdd pfet w=5 l=5
+  ad=40p pd=26u as=27p ps=16u
M1025 vdd a_690_700# A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c vdd pfet w=5 l=5
+  ad=27p pd=16u as=40p ps=26u
M1026 vdd D3 and_b2e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1027 vdd A3e_xnor_B3e A3_eq_B3_A2_eq_B2_A1_gt_B1_c vdd pfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1028 vdd D3 and_a3e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1029 A0e_xnor_B0e xor_4 gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1030 compare_A3e_nand D2 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1031 B0c compare_B0e vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1032 gnd compare_A1e A1c Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1033 and_b0e_nand B0 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1034 DEC_D2_NAND S0c DEC_AND_NODE_3 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1035 A3_eq_B3_A2_eq_B2_A1_gt_B1_c compare_A1e vdd vdd pfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1036 D3 DEC_D3_NAND vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1037 vdd D3 and_b0e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1038 and_b3e_nand B3 ander_node_8 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1039 DEC_AND_NODE_3 S1 gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1040 vdd compare_B3e_nand compare_B3e vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1041 gnd B1c A_greater_B_node_5 Gnd nfet w=5 l=5
+  ad=40p pd=26u as=27p ps=16u
M1042 and_a0e_nand A0 ander_node_4 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1043 compare_A2e_nand D2 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1044 gnd compare_A2e_nand compare_A2e Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1045 xnor_5 compare_A2e vdd vdd pfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1046 compare_node_8 B3 compare_B3e_nand Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1047 compare_node_6 B1 compare_B1e_nand Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1048 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c a_706_699# vdd vdd pfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1049 vdd A3_eq_B3_A2_gt_B2_c A3_eq_B3_A2_gt_B2 vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1050 ander_node_8 D3 gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1051 DEC_D1_NAND S1c vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1052 ander_node_4 D3 gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1053 A1_and_B1 A1_and_B1_nand vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1054 vdd A2 compare_A2e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1055 S0c S0 gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1056 A_greater_B_node_9 A2e_xnor_B2e A_greater_B_node_10 Gnd nfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1057 xnor_15 A0c gnd Gnd nfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1058 vdd S0 DEC_D1_NAND vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1059 A0e_xnor_B0e xor_4 vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1060 compare_B0e_nand D2 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1061 and_a3e and_a3e_nand gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1062 A0_and_B0 A0_and_B0_nand gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1063 gnd compare_A0e_nand compare_A0e Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1064 vdd B0 compare_B0e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1065 gnd D2 compare_node_3 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1066 gnd compare_A3e A3c Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1067 gnd A3_eq_B3_A2_eq_B2_A1_gt_B1_c A3_eq_B3_A2_eq_B2_A1_gt_B1 Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1068 S0c S0 vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1069 D3 DEC_D3_NAND gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1070 A3_eq_B3_A2_eq_B2_A1_gt_B1_c A2e_xnor_B2e vdd vdd pfet w=5 l=5
+  ad=27p pd=16u as=40p ps=26u
M1071 compare_B2e_nand D2 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1072 ander_node_10 and_b2e gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1073 gnd compare_A2e A2c Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1074 xnor_14 compare_B0e gnd Gnd nfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1075 A_compare_B_node_3 A3e_xnor_B3e A_equal_B_c Gnd nfet w=5 l=5
+  ad=27p pd=16u as=35p ps=24u
M1076 gnd compare_B0e_nand compare_B0e Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1077 A3_and_B3_nand and_a3e ander_node_9 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1078 xor_4 B0c xnor_15 Gnd nfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1079 xnor_11 compare_B1e vdd vdd pfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1080 A_equal_B_c A1e_xnor_B1e vdd vdd pfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1081 vdd B2 compare_B2e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1082 a_840_939# A_GT_B vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1083 A2_and_B2_nand and_a2e ander_node_10 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1084 A1_and_B1 A1_and_B1_nand gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1085 gnd D2 compare_node_4 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1086 A_greater_B_node_11 a_690_700# A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c Gnd nfet w=5 l=5
+  ad=27p pd=16u as=40p ps=26u
M1087 xor_2 B2c xnor_5 vdd pfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1088 vdd compare_A0e_nand compare_A0e vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1089 A_greater_B_node_6 A3e_xnor_B3e A_greater_B_node_7 Gnd nfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1090 ander_node_9 and_b3e gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1091 D0 DEC_D0_NAND gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1092 gnd A3_and_B3c A_GT_B_c Gnd nfet w=5 l=5
+  ad=40p pd=26u as=27p ps=16u
M1093 compare_node_4 A0 compare_A0e_nand Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1094 gnd compare_B2e_nand compare_B2e Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1095 vdd A3_eq_B3_A2_eq_B2_A1_gt_B1_c A3_eq_B3_A2_eq_B2_A1_gt_B1 vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1096 and_a0e and_a0e_nand vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1097 and_b3e and_b3e_nand vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1098 A_greater_B_node_5 compare_A1e A_greater_B_node_6 Gnd nfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1099 gnd compare_A1e_nand compare_A1e Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1100 vdd A3 compare_A3e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1101 A_GT_B A_GT_B_c gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1102 vdd compare_A3e A3c vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1103 vdd compare_A2e A2c vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1104 DEC_D1_NAND S1c Dec_AND_node_2 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1105 vdd compare_B0e_nand compare_B0e vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1106 vdd A3e_xnor_B3e A3_eq_B3_A2_gt_B2_c vdd pfet w=5 l=5
+  ad=40p pd=26u as=27p ps=16u
M1107 A_greater_B_node_10 a_706_699# A_greater_B_node_11 Gnd nfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1108 Dec_AND_node_2 S0 gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1109 vdd a_840_939# A_LS_B_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1110 D0 DEC_D0_NAND vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1111 compare_B1e_nand D2 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1112 xor_3 A1c xnor_11 vdd pfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1113 vdd compare_B2e_nand compare_B2e vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1114 A3_nand_B3c compare_A3e vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1115 xnor_4 compare_B3e vdd vdd pfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1116 and_b1e_nand B1 ander_node_6 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1117 xnor_13 compare_A0e vdd vdd pfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1118 gnd compare_A3e_nand compare_A3e Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1119 A1_and_B1_nand and_a1e vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1120 vdd compare_A1e_nand compare_A1e vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1121 and_a1e and_a1e_nand vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1122 xnor_8 compare_B2e vdd vdd pfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1123 xnor_12 A1c gnd Gnd nfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1124 ander_node_6 D3 gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1125 compare_node_3 A1 compare_A1e_nand Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1126 A_GT_B_c A3_and_B3c A_GT_B_node_1 vdd pfet w=5 l=5
+  ad=40p pd=26u as=27p ps=16u
M1127 A1e_xnor_B1e xor_3 vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1128 gnd A3_eq_B3_A2_eq_B2_A1_gt_B1 A_GT_B_c Gnd nfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1129 and_a0e and_a0e_nand gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1130 and_b2e and_b2e_nand vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1131 and_b3e and_b3e_nand gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1132 D1 DEC_D1_NAND vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1133 A_greater_B_node_7 A2e_xnor_B2e A3_eq_B3_A2_eq_B2_A1_gt_B1_c Gnd nfet w=5 l=5
+  ad=27p pd=16u as=35p ps=24u
M1134 gnd A3_nand_B3c A3_and_B3c Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1135 A3_and_B3 A3_and_B3_nand vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1136 B1c compare_B1e gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1137 gnd D2 compare_node_7 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1138 A_GT_B_c A3_eq_B3_A2_gt_B2 gnd Gnd nfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1139 vdd a_754_699# A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c vdd pfet w=5 l=5
+  ad=40p pd=26u as=27p ps=16u
M1140 and_b2e_nand B2 ander_node_7 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1141 vdd compare_A2e_nand compare_A2e vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1142 xnor_10 compare_B1e gnd Gnd nfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1143 and_a3e_nand A3 ander_node_1 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1144 ander_node_2 D3 gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1145 compare_node_7 B2 compare_B2e_nand Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1146 and_a2e_nand A2 ander_node_2 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1147 and_b0e and_b0e_nand vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1148 ander_node_7 D3 gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1149 gnd A0e_xnor_B0e A_compare_B_node_1 Gnd nfet w=5 l=5
+  ad=40p pd=26u as=27p ps=16u
M1150 ander_node_1 D3 gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1151 gnd compare_A0e A0c Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1152 gnd D2 compare_node_1 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1153 A3_eq_B3_A2_gt_B2_c B2c vdd vdd pfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1154 xor_1 A3c xnor_4 vdd pfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1155 and_b0e_nand B0 ander_node_5 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1156 xor_4 B0c xnor_13 vdd pfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1157 vdd A2e_xnor_B2e A_equal_B_c vdd pfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1158 vdd A3_nand_B3c A3_and_B3c vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1159 xor_2 A2c xnor_8 vdd pfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1160 DEC_D3_NAND S1 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1161 xor_3 B1c xnor_12 Gnd nfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1162 A0_and_B0_nand and_a0e vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1163 ander_node_5 D3 gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1164 xnor_16 compare_B0e vdd vdd pfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1165 gnd D2 compare_node_2 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1166 xnor_3 A3c gnd Gnd nfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1167 and_a1e and_a1e_nand gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1168 vdd S0 DEC_D3_NAND vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1169 A_GT_B_node_2 A3_eq_B3_A2_eq_B2_A1_gt_B1 A_GT_B_node_3 vdd pfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1170 gnd A3e_xnor_B3e A_greater_B_node_2 Gnd nfet w=5 l=5
+  ad=40p pd=26u as=27p ps=16u
M1171 vdd and_b0e A0_and_B0_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1172 A1e_xnor_B1e xor_3 gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1173 D2 DEC_D2_NAND vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1174 DEC_D2_NAND S0c vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1175 compare_B3e_nand D2 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1176 compare_node_2 A2 compare_A2e_nand Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1177 and_b2e and_b2e_nand gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1178 D1 DEC_D1_NAND gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1179 A_LS_B_node_1 a_840_939# A_LS_B_nand Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1180 and_b3e_nand B3 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1181 vdd compare_A0e A0c vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1182 vdd S1 DEC_D2_NAND vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1183 A3_and_B3 A3_and_B3_nand gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1184 xor_3 compare_A1e xnor_10 Gnd nfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1185 A_GT_B_node_1 A3_eq_B3_A2_gt_B2 A_GT_B_node_2 vdd pfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1186 gnd compare_A3e A_greater_B_node_1 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1187 xnor_2 compare_B3e gnd Gnd nfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1188 vdd D3 and_b3e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1189 and_b1e and_b1e_nand vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1190 gnd D2 compare_node_5 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1191 vdd B1 compare_B1e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1192 vdd B3c A3_nand_B3c vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1193 xnor_6 compare_B2e gnd Gnd nfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1194 A1_and_B1_nand and_a1e ander_node_11 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1195 and_b0e and_b0e_nand gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1196 compare_node_5 B0 compare_B0e_nand Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1197 A_GT_B_c A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 gnd Gnd nfet w=5 l=5
+  ad=27p pd=16u as=40p ps=26u
M1198 xor_4 compare_A0e xnor_14 Gnd nfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1199 DEC_D0_NAND S0c vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1200 A2_and_B2 A2_and_B2_nand vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1201 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c A3e_xnor_B3e vdd vdd pfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1202 xor_1 B3c xnor_3 Gnd nfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1203 vdd and_b1e A1_and_B1_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1204 xnor_9 compare_A1e vdd vdd pfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1205 gnd a_754_699# A_greater_B_node_8 Gnd nfet w=5 l=5
+  ad=40p pd=26u as=27p ps=16u
M1206 vdd S1c DEC_D0_NAND vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1207 and_a1e_nand A1 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1208 vdd and_b2e A2_and_B2_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1209 compare_A1e_nand D2 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1210 A3e_xnor_B3e xor_1 gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1211 A3_and_B3_nand and_a3e vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1212 A_GT_B A_GT_B_c vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1213 gnd A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1214 A2_and_B2_nand and_a2e vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1215 D2 DEC_D2_NAND gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1216 A_compare_B_node_1 A1e_xnor_B1e A_compare_B_node_2 Gnd nfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1217 gnd compare_B1e_nand compare_B1e Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1218 A_LS_B_nand A_equal_B_c vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1219 vdd D3 and_a1e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1220 S1c S1 gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1221 vdd and_b3e A3_and_B3_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1222 gnd A_equal_B_c A_equal_B Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1223 vdd compare_A2e A3_eq_B3_A2_gt_B2_c vdd pfet w=5 l=5
+  ad=27p pd=16u as=40p ps=26u
M1224 xor_1 compare_A3e xnor_2 Gnd nfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1225 A_greater_B_node_2 B2c A_greater_B_node_3 Gnd nfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1226 and_a2e and_a2e_nand vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1227 A_equal_B_c A3e_xnor_B3e vdd vdd pfet w=5 l=5
+  ad=27p pd=16u as=40p ps=26u
M1228 and_b1e and_b1e_nand gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1229 DEC_D3_NAND S1 DEC_AND_NODE_4 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1230 compare_A0e_nand D2 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1231 A2e_xnor_B2e xor_2 gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1232 gnd A_LS_B_nand A_LS_B Gnd nfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1233 A0_and_B0_nand and_a0e ander_node_12 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1234 vdd compare_A3e_nand compare_A3e vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1235 DEC_AND_NODE_4 S0 gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1236 A_GT_B_node_3 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 vdd vdd pfet w=5 l=5
+  ad=27p pd=16u as=40p ps=26u
M1237 vdd A0 compare_A0e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1238 xor_2 compare_A2e xnor_6 Gnd nfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1239 compare_node_1 A3 compare_A3e_nand Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1240 vdd A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1241 ander_node_12 and_b0e gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1242 gnd D2 compare_node_8 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1243 xnor_7 A2c gnd Gnd nfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1244 vdd compare_B1e_nand compare_B1e vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1245 A2_and_B2 A2_and_B2_nand gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1246 xor_3 B1c xnor_9 vdd pfet w=5 l=5
+  ad=40p pd=26u as=32p ps=18u
M1247 S1c S1 vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1248 vdd A_equal_B_c A_equal_B vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1249 vdd B1c A3_eq_B3_A2_eq_B2_A1_gt_B1_c vdd pfet w=5 l=5
+  ad=40p pd=26u as=27p ps=16u
M1250 xnor_1 compare_A3e vdd vdd pfet w=5 l=5
+  ad=32p pd=18u as=40p ps=26u
M1251 and_a0e_nand A0 vdd vdd pfet w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1252 B1c compare_B1e vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1253 gnd D2 compare_node_6 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1254 A_greater_B_node_1 B3c A3_nand_B3c Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1255 a_840_939# A_GT_B gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1256 vdd B3 compare_B3e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1257 A3e_xnor_B3e xor_1 vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1258 vdd D3 and_a0e_nand vdd pfet w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1259 A2e_xnor_B2e xor_2 vdd vdd pfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1260 vdd A_LS_B_nand A_LS_B vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1261 vdd A2e_xnor_B2e A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c vdd pfet w=5 l=5
+  ad=27p pd=16u as=27p ps=16u
M1262 B3c compare_B3e gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1263 vdd compare_A1e A1c vdd pfet w=5 l=5
+  ad=35p pd=24u as=40p ps=26u
M1264 and_a2e and_a2e_nand gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1265 DEC_D0_NAND S0c Dec_AND_node_1 Gnd nfet w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1266 B2c compare_B2e gnd Gnd nfet w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1267 ander_node_11 and_b1e gnd Gnd nfet w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
C0 A3e_xnor_B3e B3c 0.051034f
C1 ander_node_8 D3 0.089107f
C2 xor_4 vdd 0.515131f
C3 gnd A2e_xnor_B2e 0.071179f
C4 A3_eq_B3_A2_eq_B2_A1_gt_B1 B1c 0.79062f
C5 gnd and_b3e 0.081083f
C6 A3_eq_B3_A2_gt_B2 vdd 0.126896f
C7 gnd Dec_AND_node_1 0.07683f
C8 D2 compare_node_2 0.089107f
C9 A0e_xnor_B0e xor_4 0.036f
C10 and_b1e D3 0.007976f
C11 and_a2e A0 0.010567f
C12 and_a1e_nand D3 0.015311f
C13 xor_4 xnor_15 1.47e-19
C14 B0 compare_B1e 0.013715f
C15 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 B1c 0.08784f
C16 S0c DEC_D2_NAND 0.006448f
C17 A2e_xnor_B2e A_equal_B_c 0.017948f
C18 and_a2e vdd 0.135377f
C19 ander_node_1 A3 0.088221f
C20 A2e_xnor_B2e B3c 0.023722f
C21 A2e_xnor_B2e A3e_xnor_B3e 0.32451f
C22 compare_A3e compare_A3e_nand 0.030251f
C23 a_754_699# compare_A0e 0.012143f
C24 gnd A1_and_B1 0.051616f
C25 A0_and_B0_nand A0_and_B0 0.030251f
C26 and_b0e ander_node_12 0.089107f
C27 and_a2e ander_node_10 0.088221f
C28 S1c Dec_AND_node_2 0.088221f
C29 B2c compare_A3e 0.090491f
C30 and_b2e_nand D3 0.015311f
C31 a_754_699# vdd 0.075131f
C32 gnd B3 0.012704f
C33 A_GT_B_c A3_and_B3c 0.027212f
C34 A0_and_B0 vdd 0.040884f
C35 and_a1e and_a0e 0.012215f
C36 and_b2e and_b0e 0.01764f
C37 ander_node_7 D3 0.089107f
C38 gnd A0_and_B0_nand 0.148342f
C39 B2 vdd 0.151575f
C40 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 A1e_xnor_B1e 0.056906f
C41 gnd compare_A0e 0.218845f
C42 B1c compare_B1e 0.030251f
C43 and_a3e and_a2e 0.029024f
C44 gnd A0 0.131974f
C45 compare_A0e compare_B3e 0.011781f
C46 gnd a_690_700# 0.015532f
C47 gnd xnor_3 1.47e-19
C48 gnd vdd 0.286842f
C49 compare_A2e_nand vdd 0.094003f
C50 compare_B3e vdd 0.162042f
C51 S1c DEC_D1_NAND 0.006448f
C52 compare_B1e_nand compare_B1e 0.030251f
C53 A3 D3 0.112603f
C54 gnd A0e_xnor_B0e 0.142939f
C55 compare_A2e compare_B2e 0.03971f
C56 a_706_699# vdd 0.075131f
C57 gnd xnor_15 1.47e-19
C58 gnd ander_node_10 0.07683f
C59 compare_A3e A2 0.218758f
C60 A3_eq_B3_A2_gt_B2 A3_and_B3c 0.016979f
C61 and_a1e ander_node_11 0.088221f
C62 vdd A_equal_B_c 0.328347f
C63 D2 B2 0.007976f
C64 compare_B1e_nand compare_node_6 0.085282f
C65 ander_node_4 A0 0.08968f
C66 compare_A3e A3_nand_B3c 0.015311f
C67 B0c compare_A0e 0.021235f
C68 A0e_xnor_B0e A_equal_B_c 0.003222f
C69 B3c vdd 0.46262f
C70 A3e_xnor_B3e vdd 0.989055f
C71 gnd A3_and_B3_nand 0.148342f
C72 gnd compare_B3e_nand 0.148342f
C73 D2 gnd 0.334121f
C74 and_a2e_nand and_a2e 0.030251f
C75 D2 compare_node_7 0.089107f
C76 D2 compare_A2e_nand 0.015311f
C77 compare_A1e A1c 0.038705f
C78 compare_B3e_nand compare_B3e 0.030251f
C79 D2 compare_B3e 0.005588f
C80 B0c vdd 0.212299f
C81 gnd compare_node_8 0.07683f
C82 gnd and_a3e 0.051616f
C83 gnd A_greater_B_node_2 6.22e-20
C84 D0 vdd 0.040884f
C85 and_a2e A1 0.077299f
C86 and_b2e_nand ander_node_7 0.085282f
C87 gnd A3_eq_B3_A2_eq_B2_A1_gt_B1_c 0.058859f
C88 A2e_xnor_B2e vdd 1.24529f
C89 gnd compare_node_1 0.07683f
C90 and_b3e vdd 0.11701f
C91 B0 and_b2e 0.007976f
C92 DEC_D1_NAND D1 0.030251f
C93 gnd DEC_D2_NAND 0.157853f
C94 S1 DEC_AND_NODE_4 0.088221f
C95 gnd A2_and_B2 0.051616f
C96 and_a0e ander_node_12 0.088221f
C97 and_b0e_nand gnd 0.148342f
C98 a_840_939# A_LS_B_nand 0.006448f
C99 S1c S1 0.030251f
C100 ander_node_3 D3 0.089107f
C101 A3_eq_B3_A2_gt_B2_c compare_A2e 0.0242f
C102 A3e_xnor_B3e A3_eq_B3_A2_eq_B2_A1_gt_B1_c 0.017948f
C103 A_LS_B_node_1 A_LS_B_nand 0.085282f
C104 gnd A3_and_B3c 0.136884f
C105 A1_and_B1 vdd 0.040884f
C106 gnd and_a2e_nand 0.148342f
C107 and_b3e A3_and_B3_nand 0.015311f
C108 and_a1e_nand and_a1e 0.030251f
C109 ander_node_5 gnd 0.07683f
C110 compare_B0e compare_B2e 0.008162f
C111 DEC_AND_NODE_4 S0 0.089107f
C112 A_LS_B A_LS_B_nand 0.030251f
C113 A3_eq_B3_A2_gt_B2 B2c 0.001885f
C114 B3 vdd 0.151897f
C115 gnd xnor_7 1.47e-19
C116 S1c S0 0.07308f
C117 gnd A1 0.076253f
C118 A3_and_B3c B3c 0.008592f
C119 A2e_xnor_B2e A3_eq_B3_A2_eq_B2_A1_gt_B1_c 0.029291f
C120 A0_and_B0_nand vdd 0.094003f
C121 compare_A0e vdd 0.176676f
C122 ander_node_1 and_a3e_nand 0.085282f
C123 and_a1e_nand ander_node_3 0.085282f
C124 compare_node_2 A2 0.088221f
C125 A0 vdd 0.197884f
C126 and_b3e_nand gnd 0.148342f
C127 compare_B0e compare_B1e 0.014402f
C128 a_690_700# vdd 0.075131f
C129 A1_and_B1_nand ander_node_11 0.085282f
C130 compare_A3e A_greater_B_node_1 0.089107f
C131 compare_B3e_nand B3 0.006448f
C132 D2 B3 0.016016f
C133 gnd compare_B0e_nand 0.148342f
C134 S1c DEC_D0_NAND 0.015311f
C135 compare_A3e compare_A2e 0.182612f
C136 A0e_xnor_B0e vdd 0.139586f
C137 compare_node_8 B3 0.088221f
C138 gnd and_b0e 0.113067f
C139 A2c gnd 1.43721f
C140 and_a0e_nand and_a0e 0.030251f
C141 and_b2e A2_and_B2_nand 0.015311f
C142 compare_B1e compare_B2e 0.015731f
C143 compare_A1e xor_3 0.008861f
C144 gnd A_equal_B 0.051616f
C145 gnd compare_A3e_nand 0.148342f
C146 A3_and_B3_nand vdd 0.094003f
C147 D2 vdd 0.673071f
C148 compare_A1e_nand compare_node_3 0.085282f
C149 compare_B3e_nand vdd 0.094003f
C150 and_b2e D3 0.00917f
C151 and_a3e A0 0.013687f
C152 gnd B2c 0.174287f
C153 S1 DEC_AND_NODE_3 0.089107f
C154 and_a3e vdd 0.14109f
C155 A_equal_B A_equal_B_c 0.030251f
C156 B2c compare_B3e 0.020796f
C157 compare_B1e_nand B1 0.006448f
C158 and_b3e_nand and_b3e 0.030251f
C159 D3 and_a3e_nand 0.015311f
C160 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c a_754_699# 0.003222f
C161 gnd A1c 1.43721f
C162 S1 DEC_D3_NAND 0.006448f
C163 A3_eq_B3_A2_eq_B2_A1_gt_B1_c vdd 0.227022f
C164 gnd A3_and_B3 0.051616f
C165 D2 compare_B3e_nand 0.015311f
C166 S0c S1 0.511187f
C167 compare_A1e compare_A2e 0.030403f
C168 A3e_xnor_B3e B2c 0.293828f
C169 B2c B3c 0.07507f
C170 A_LS_B_node_1 a_840_939# 0.088221f
C171 DEC_D2_NAND vdd 0.094003f
C172 DEC_D3_NAND D3 0.030251f
C173 and_b1e A1_and_B1_nand 0.015311f
C174 A2_and_B2 vdd 0.040884f
C175 A2c A2e_xnor_B2e 0.041238f
C176 gnd Dec_AND_node_2 0.077312f
C177 and_b2e and_b1e 0.010402f
C178 and_b3e and_b0e 0.01764f
C179 and_a2e and_a0e 0.008592f
C180 and_a3e A3_and_B3_nand 0.006448f
C181 D2 compare_node_8 0.089107f
C182 compare_B3e_nand compare_node_8 0.085282f
C183 B1 D3 0.0056f
C184 and_b0e_nand vdd 0.094003f
C185 DEC_D3_NAND S0 0.015311f
C186 gnd A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c 0.058859f
C187 gnd compare_node_4 0.07683f
C188 A3_and_B3c vdd 0.126682f
C189 D2 compare_node_1 0.089107f
C190 S0c S0 0.043542f
C191 and_a2e_nand vdd 0.094003f
C192 gnd A2 0.102362f
C193 and_a0e_nand D3 0.015311f
C194 and_b3e_nand B3 0.006448f
C195 compare_A2e_nand A2 0.006448f
C196 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c a_706_699# 0.020823f
C197 gnd A3_nand_B3c 0.162217f
C198 A2e_xnor_B2e B2c 0.004638f
C199 D2 DEC_D2_NAND 0.030251f
C200 compare_B0e A0c 0.014332f
C201 gnd ander_node_2 0.07683f
C202 A1 vdd 0.21183f
C203 B0 gnd 0.00543f
C204 and_b2e_nand and_b2e 0.030251f
C205 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c A3e_xnor_B3e 0.017948f
C206 B0 compare_B3e 0.004394f
C207 gnd DEC_D1_NAND 0.159401f
C208 S0c DEC_D0_NAND 0.006448f
C209 and_b3e_nand vdd 0.094003f
C210 compare_A3e A3c 0.040434f
C211 B3c A3_nand_B3c 0.006448f
C212 A_GT_B a_840_939# 0.030251f
C213 and_b1e_nand D3 0.015311f
C214 gnd and_a0e 0.083816f
C215 and_b0e A0_and_B0_nand 0.015311f
C216 and_a2e A2_and_B2_nand 0.006448f
C217 xor_2 gnd 0.127657f
C218 gnd compare_A0e_nand 0.148342f
C219 compare_B0e_nand vdd 0.094003f
C220 xor_3 xnor_12 1.47e-19
C221 ander_node_6 D3 0.089107f
C222 A2e_xnor_B2e A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c 0.017948f
C223 gnd ander_node_1 0.07683f
C224 and_b0e vdd 0.116913f
C225 A2c vdd 0.146829f
C226 and_a3e A1 0.010584f
C227 gnd B1c 0.630143f
C228 A_equal_B vdd 0.04098f
C229 compare_A3e_nand vdd 0.094003f
C230 and_b1e_nand and_b1e 0.030251f
C231 D2 compare_B0e_nand 0.015311f
C232 B0 and_b3e 0.005588f
C233 and_b0e_nand ander_node_5 0.085282f
C234 A3 and_a3e_nand 0.006448f
C235 gnd xor_3 0.127657f
C236 compare_A1e compare_B2e 0.012373f
C237 B2c vdd 0.429881f
C238 gnd ander_node_11 0.07683f
C239 A_GT_B_c A3_eq_B3_A2_eq_B2_A1_gt_B1 0.018351f
C240 gnd compare_B1e_nand 0.148342f
C241 B1c B3c 0.017541f
C242 A3e_xnor_B3e B1c 0.036396f
C243 A1c vdd 0.146829f
C244 B1 compare_B2e 0.010094f
C245 A_GT_B_c A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 0.003625f
C246 gnd A2_and_B2_nand 0.148342f
C247 xor_2 A2e_xnor_B2e 0.036f
C248 A3_and_B3 vdd 0.040884f
C249 and_a1e A1_and_B1_nand 0.006448f
C250 gnd S1 0.131827f
C251 compare_B2e_nand compare_B2e 0.030251f
C252 D2 compare_A3e_nand 0.015311f
C253 B2 D3 0.006732f
C254 A0e_xnor_B0e A1c 0.03623f
C255 gnd A1e_xnor_B1e 0.233988f
C256 compare_A1e compare_B1e 0.036091f
C257 gnd D3 0.313918f
C258 gnd A_greater_B_node_1 0.077137f
C259 compare_node_4 A0 0.088221f
C260 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c a_690_700# 0.029281f
C261 A2e_xnor_B2e B1c 0.005883f
C262 gnd compare_A2e 0.252662f
C263 compare_A2e compare_A2e_nand 0.030251f
C264 gnd S0 0.110102f
C265 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c vdd 0.264836f
C266 compare_A3e_nand compare_node_1 0.085282f
C267 A1e_xnor_B1e A_equal_B_c 0.017948f
C268 compare_A2e compare_B3e 0.02951f
C269 A3_and_B3_nand A3_and_B3 0.030251f
C270 A3_eq_B3_A2_eq_B2_A1_gt_B1 A3_eq_B3_A2_gt_B2 0.063504f
C271 A2 vdd 0.207071f
C272 and_b0e_nand and_b0e 0.030251f
C273 B3c A1e_xnor_B1e 0.093078f
C274 A3e_xnor_B3e A1e_xnor_B1e 0.018378f
C275 A3_nand_B3c vdd 0.094003f
C276 B3c A_greater_B_node_1 0.088221f
C277 compare_node_6 B1 0.088221f
C278 gnd compare_node_5 0.07683f
C279 ander_node_8 gnd 0.07683f
C280 ander_node_4 D3 0.089107f
C281 B0 vdd 0.151575f
C282 xor_1 A3c 0.03574f
C283 gnd A_LS_B_nand 0.148342f
C284 gnd and_b1e 0.102119f
C285 and_a0e A0_and_B0_nand 0.006448f
C286 gnd and_a1e_nand 0.148342f
C287 DEC_D0_NAND gnd 0.145266f
C288 D2 compare_node_4 0.089107f
C289 compare_A2e B0c 0.030873f
C290 compare_A0e_nand compare_A0e 0.030251f
C291 DEC_D1_NAND vdd 0.094035f
C292 compare_A0e_nand A0 0.006448f
C293 A_LS_B_nand A_equal_B_c 0.015311f
C294 A2e_xnor_B2e A1e_xnor_B1e 0.012877f
C295 gnd compare_node_3 0.07683f
C296 and_a0e vdd 0.136432f
C297 xor_2 vdd 0.452209f
C298 DEC_D3_NAND DEC_AND_NODE_4 0.085282f
C299 compare_A0e_nand vdd 0.094003f
C300 and_b3e D3 0.006732f
C301 and_a3e A2 0.164509f
C302 and_b2e_nand B2 0.006448f
C303 B0 D2 0.004411f
C304 compare_A1e compare_A1e_nand 0.030251f
C305 ander_node_7 B2 0.088221f
C306 and_b2e_nand gnd 0.148342f
C307 S0c S1c 0.015985f
C308 B1c vdd 0.644935f
C309 gnd A3_eq_B3_A2_eq_B2_A1_gt_B1 0.117028f
C310 ander_node_7 gnd 0.07683f
C311 gnd compare_B0e 0.702733f
C312 DEC_D0_NAND D0 0.030251f
C313 D2 compare_A0e_nand 0.015311f
C314 compare_A1e compare_A3e 0.012373f
C315 compare_B0e compare_B3e 0.008162f
C316 xor_3 vdd 0.531725f
C317 A_GT_B_c A_GT_B 0.030251f
C318 gnd A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 0.117028f
C319 and_b3e and_b1e 0.010402f
C320 and_a3e and_a0e 0.012211f
C321 and_a2e and_a1e 0.010267f
C322 B3 D3 0.004542f
C323 DEC_D0_NAND Dec_AND_node_1 0.085282f
C324 compare_B1e_nand vdd 0.094003f
C325 and_a2e_nand A2 0.006448f
C326 B0 and_b0e_nand 0.006448f
C327 A3_and_B3c A3_nand_B3c 0.030251f
C328 A3_eq_B3_A2_eq_B2_A1_gt_B1 B3c 0.017618f
C329 A3_eq_B3_A2_gt_B2 A3_eq_B3_A2_gt_B2_c 0.030251f
C330 A3_eq_B3_A2_eq_B2_A1_gt_B1 A3e_xnor_B3e 0.035581f
C331 gnd compare_B2e 0.281f
C332 A2_and_B2_nand vdd 0.094003f
C333 S1 vdd 0.201098f
C334 gnd A3 0.010267f
C335 and_a2e_nand ander_node_2 0.085282f
C336 compare_B2e compare_B3e 0.004394f
C337 A2 A1 0.02262f
C338 B0 ander_node_5 0.088221f
C339 gnd A3c 1.43721f
C340 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 A3e_xnor_B3e 0.034381f
C341 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 B3c 0.029257f
C342 a_690_700# A1e_xnor_B1e 0.006476f
C343 compare_B0e B0c 0.030251f
C344 compare_A2e compare_A0e 0.036913f
C345 A1e_xnor_B1e vdd 0.208204f
C346 A3c compare_B3e 0.014332f
C347 A2_and_B2_nand ander_node_10 0.085282f
C348 compare_A2e A0 0.03114f
C349 ander_node_8 B3 0.088221f
C350 D3 vdd 0.659484f
C351 D2 compare_B1e_nand 0.015311f
C352 B1c A3_eq_B3_A2_eq_B2_A1_gt_B1_c 0.003222f
C353 A1e_xnor_B1e A0e_xnor_B0e 0.229516f
C354 compare_A2e vdd 0.282244f
C355 S0 vdd 0.202099f
C356 and_b2e B1 0.010094f
C357 A3_eq_B3_A2_eq_B2_A1_gt_B1 A2e_xnor_B2e 0.020477f
C358 gnd compare_B1e 0.28163f
C359 xor_1 compare_A3e 0.008861f
C360 A3e_xnor_B3e A3c 0.041238f
C361 B0c compare_B2e 0.021297f
C362 compare_B1e compare_B3e 0.004394f
C363 gnd a_840_939# 0.060377f
C364 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 A2e_xnor_B2e 0.052742f
C365 A_LS_B_node_1 gnd 0.07683f
C366 gnd and_a1e 0.084316f
C367 gnd compare_node_6 0.07683f
C368 xor_2 xnor_7 1.47e-19
C369 D2 D3 0.010267f
C370 A_LS_B_nand vdd 0.094003f
C371 B0 compare_B0e_nand 0.006448f
C372 A_LS_B gnd 0.051616f
C373 S0c DEC_AND_NODE_3 0.088221f
C374 A_LS_B_node_1 A_equal_B_c 0.089107f
C375 and_b1e vdd 0.11701f
C376 and_a1e_nand vdd 0.094003f
C377 xor_4 A0c 0.03574f
C378 DEC_D0_NAND vdd 0.094023f
C379 and_a3e D3 1.7e-20
C380 gnd A3_eq_B3_A2_gt_B2_c 0.139896f
C381 compare_B1e B0c 0.020681f
C382 S1 DEC_D2_NAND 0.015311f
C383 A2_and_B2_nand A2_and_B2 0.030251f
C384 gnd ander_node_3 0.07683f
C385 D2 compare_node_5 0.089107f
C386 gnd DEC_AND_NODE_4 0.077062f
C387 S1c gnd 0.055406f
C388 xor_2 A2c 0.03574f
C389 compare_B0e compare_A0e 0.142568f
C390 and_b2e_nand vdd 0.094003f
C391 A3e_xnor_B3e A3_eq_B3_A2_gt_B2_c 0.003222f
C392 and_b0e_nand D3 0.015311f
C393 gnd A_GT_B 0.113911f
C394 gnd compare_A1e_nand 0.148342f
C395 A3_eq_B3_A2_eq_B2_A1_gt_B1 vdd 0.162801f
C396 D2 compare_node_3 0.089107f
C397 compare_B0e vdd 0.162042f
C398 and_a2e_nand D3 0.015311f
C399 ander_node_5 D3 0.089107f
C400 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 vdd 0.205943f
C401 xor_2 B2c 0.075488f
C402 compare_A0e compare_B2e 0.014064f
C403 and_b1e_nand B1 0.006448f
C404 gnd compare_A3e 0.156193f
C405 compare_B2e vdd 0.162042f
C406 compare_A3e compare_B3e 0.046926f
C407 compare_A2e A1 0.137799f
C408 ander_node_6 B1 0.088221f
C409 A3 vdd 0.226675f
C410 ander_node_2 A2 0.091719f
C411 DEC_D1_NAND Dec_AND_node_2 0.085282f
C412 gnd A0c 1.43721f
C413 B1c B2c 0.068709f
C414 and_b3e_nand D3 0.015311f
C415 A3c vdd 0.146105f
C416 gnd ander_node_12 0.07683f
C417 A_GT_B_c A3_eq_B3_A2_gt_B2 0.018351f
C418 gnd D1 0.051616f
C419 compare_B1e compare_A0e 0.020796f
C420 S1c Dec_AND_node_1 0.089107f
C421 A3_eq_B3_A2_eq_B2_A1_gt_B1 A3_eq_B3_A2_eq_B2_A1_gt_B1_c 0.030251f
C422 gnd and_b2e 0.114913f
C423 gnd A1_and_B1_nand 0.148342f
C424 D2 compare_B2e 0.004394f
C425 compare_A0e_nand compare_node_4 0.085282f
C426 compare_B1e vdd 0.162042f
C427 compare_A3e B0c 0.015831f
C428 and_a1e A0 0.006955f
C429 xor_3 A1c 0.03574f
C430 and_a1e_nand A1 0.006448f
C431 a_840_939# vdd 0.275571f
C432 and_b3e_nand ander_node_8 0.085282f
C433 A2c compare_A2e 0.038705f
C434 and_a1e vdd 0.144029f
C435 gnd and_a3e_nand 0.148342f
C436 compare_node_3 A1 0.088951f
C437 and_b1e_nand ander_node_6 0.085282f
C438 compare_B0e_nand compare_node_5 0.085282f
C439 gnd DEC_AND_NODE_3 0.077196f
C440 gnd compare_A1e 0.29778f
C441 B2c A1e_xnor_B1e 0.127099f
C442 A_LS_B vdd 0.04098f
C443 gnd ander_node_9 0.07683f
C444 compare_A1e compare_B3e 0.026206f
C445 compare_B2e_nand B2 0.006448f
C446 compare_node_1 A3 0.088221f
C447 D2 compare_B1e 0.004394f
C448 gnd DEC_D3_NAND 0.157853f
C449 A1e_xnor_B1e A1c 0.049486f
C450 A3_eq_B3_A2_gt_B2_c vdd 0.188033f
C451 gnd B1 0.00875f
C452 and_b1e and_b0e 0.01764f
C453 S0c gnd 0.051616f
C454 gnd compare_B2e_nand 0.148342f
C455 B1 compare_B3e 0.007976f
C456 D2 compare_node_6 0.089107f
C457 compare_B2e_nand compare_node_7 0.085282f
C458 gnd A_GT_B_c 0.317056f
C459 gnd and_a0e_nand 0.148342f
C460 and_a3e and_a1e 0.053894f
C461 and_b3e and_b2e 0.012211f
C462 gnd A_greater_B_node_3 6.22e-20
C463 compare_A1e B0c 0.015248f
C464 S1c vdd 0.19269f
C465 gnd compare_node_2 0.07683f
C466 A_GT_B vdd 0.090595f
C467 Dec_AND_node_2 S0 0.089107f
C468 compare_A2e_nand compare_node_2 0.085282f
C469 compare_A1e_nand vdd 0.094003f
C470 compare_B0e_nand compare_B0e 0.030251f
C471 gnd xor_1 0.127657f
C472 compare_A3e compare_A0e 0.036236f
C473 A3_nand_B3c A_greater_B_node_1 0.085282f
C474 and_b3e ander_node_9 0.089107f
C475 compare_A3e A0 0.029337f
C476 A1_and_B1_nand A1_and_B1 0.030251f
C477 and_a0e_nand ander_node_4 0.085282f
C478 and_b1e_nand gnd 0.148342f
C479 ander_node_2 D3 0.089107f
C480 gnd xor_4 0.127657f
C481 A0c compare_A0e 0.038705f
C482 B0 D3 0.008116f
C483 compare_A3e vdd 0.284455f
C484 and_b3e B1 0.00709f
C485 A0_and_B0_nand ander_node_12 0.085282f
C486 gnd A3_eq_B3_A2_gt_B2 0.119903f
C487 ander_node_6 gnd 0.07683f
C488 D2 compare_A1e_nand 0.015311f
C489 S0c Dec_AND_node_1 0.088221f
C490 B3c xor_1 0.075488f
C491 B1c xor_3 0.075488f
C492 A3e_xnor_B3e xor_1 0.039012f
C493 A0c vdd 0.146829f
C494 A3_eq_B3_A2_eq_B2_A1_gt_B1 B2c 0.142748f
C495 gnd and_a2e 0.095887f
C496 DEC_D1_NAND S0 0.015311f
C497 A2c compare_B2e 0.014332f
C498 D1 vdd 0.04098f
C499 A0e_xnor_B0e A0c 0.041238f
C500 B0 compare_node_5 0.088221f
C501 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 B2c 0.11379f
C502 A3_eq_B3_A2_gt_B2 B3c 0.00709f
C503 A3_eq_B3_A2_gt_B2 A3e_xnor_B3e 0.031799f
C504 xor_2 compare_A2e 0.008861f
C505 A1_and_B1_nand vdd 0.094003f
C506 and_b2e vdd 0.11701f
C507 B0c xor_4 0.075488f
C508 ander_node_1 D3 0.089107f
C509 compare_A3e_nand A3 0.006448f
C510 B0 and_b1e 0.006782f
C511 gnd xnor_12 1.47e-19
C512 gnd a_754_699# 0.018955f
C513 compare_A1e compare_A0e 0.016585f
C514 B1c A1e_xnor_B1e 0.011342f
C515 B2c compare_B2e 0.030251f
C516 gnd A0_and_B0 0.051616f
C517 compare_A1e A0 0.260485f
C518 and_b2e ander_node_10 0.089107f
C519 and_a3e_nand vdd 0.094003f
C520 ander_node_3 A1 0.09041f
C521 B1c compare_A2e 0.016406f
C522 A1e_xnor_B1e xor_3 0.055608f
C523 compare_A1e vdd 0.265389f
C524 gnd B2 0.020143f
C525 compare_node_7 B2 0.088221f
C526 and_b1e and_a0e 4.19e-21
C527 B2 compare_B3e 0.007976f
C528 DEC_D3_NAND vdd 0.094059f
C529 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c 0.030251f
C530 B1 vdd 0.151575f
C531 gnd compare_node_7 0.07683f
C532 gnd compare_A2e_nand 0.148342f
C533 S0c vdd 0.230788f
C534 compare_B2e_nand vdd 0.094003f
C535 gnd compare_B3e 0.306994f
C536 and_a0e_nand A0 0.006448f
C537 compare_A1e_nand A1 0.006448f
C538 gnd a_706_699# 0.015532f
C539 D2 compare_A1e 1.7e-20
C540 compare_B1e A1c 0.014332f
C541 gnd A_equal_B_c 0.148523f
C542 A_GT_B_c vdd 0.070745f
C543 S1 S0 0.028532f
C544 and_a0e_nand vdd 0.094003f
C545 A3_and_B3_nand ander_node_9 0.085282f
C546 and_a3e and_a3e_nand 0.030251f
C547 gnd B3c 0.088039f
C548 gnd A3e_xnor_B3e 0.089328f
C549 gnd ander_node_4 0.07683f
C550 D2 B1 0.007988f
C551 and_a3e ander_node_9 0.088221f
C552 compare_A3e A1 0.025755f
C553 B3c compare_B3e 0.030251f
C554 and_b1e ander_node_11 0.089107f
C555 D2 compare_B2e_nand 0.015311f
C556 B0 compare_B2e 0.004394f
C557 xor_1 xnor_3 1.47e-19
C558 gnd B0c 0.689019f
C559 B2c A3_eq_B3_A2_gt_B2_c 0.020823f
C560 A3_eq_B3_A2_eq_B2_A1_gt_B1_c compare_A1e 0.017948f
C561 xor_4 compare_A0e 0.008861f
C562 xor_1 vdd 0.410409f
C563 A3e_xnor_B3e A_equal_B_c 0.029291f
C564 B0c compare_B3e 0.245979f
C565 and_b3e B2 0.105897f
C566 D0 gnd 0.051616f
C567 a_706_699# B0c 0.009511f
C568 and_b1e_nand vdd 0.094003f
C569 DEC_D2_NAND DEC_AND_NODE_3 0.085282f
C570 A0c 0 1.68244f **FLOATING
C571 xor_4 0 1.62527f **FLOATING
C572 B0c 0 3.62443f **FLOATING
C573 DEC_AND_NODE_4 0 0.248064f **FLOATING
C574 DEC_D3_NAND 0 0.516966f **FLOATING
C575 DEC_AND_NODE_3 0 0.248064f **FLOATING
C576 DEC_D2_NAND 0 0.52029f **FLOATING
C577 A1c 0 1.67561f **FLOATING
C578 xor_3 0 1.78086f **FLOATING
C579 A0e_xnor_B0e 0 2.34631f **FLOATING
C580 A1e_xnor_B1e 0 10.189f **FLOATING
C581 compare_node_8 0 0.248064f **FLOATING
C582 A_equal_B 0 0.088325f **FLOATING
C583 compare_node_7 0 0.248064f **FLOATING
C584 compare_node_6 0 0.248064f **FLOATING
C585 Dec_AND_node_2 0 0.248064f **FLOATING
C586 S1 0 2.76414f **FLOATING
C587 compare_B3e_nand 0 0.52029f **FLOATING
C588 compare_B2e_nand 0 0.52029f **FLOATING
C589 compare_node_5 0 0.248064f **FLOATING
C590 compare_B1e 0 11.4538f **FLOATING
C591 D1 0 0.104663f **FLOATING
C592 compare_B1e_nand 0 0.52029f **FLOATING
C593 compare_B0e 0 7.35184f **FLOATING
C594 compare_B0e_nand 0 0.52029f **FLOATING
C595 DEC_D1_NAND 0 0.513722f **FLOATING
C596 S0 0 7.9098f **FLOATING
C597 compare_node_1 0 0.248064f **FLOATING
C598 compare_node_2 0 0.248064f **FLOATING
C599 compare_node_3 0 0.248064f **FLOATING
C600 compare_node_4 0 0.248064f **FLOATING
C601 compare_B2e 0 13.3011f **FLOATING
C602 compare_A3e_nand 0 0.52029f **FLOATING
C603 compare_A2e_nand 0 0.52029f **FLOATING
C604 compare_A0e 0 13.6565f **FLOATING
C605 Dec_AND_node_1 0 0.248064f **FLOATING
C606 compare_A1e_nand 0 0.52029f **FLOATING
C607 compare_A0e_nand 0 0.52029f **FLOATING
C608 D0 0 0.395495f **FLOATING
C609 D2 0 28.4675f **FLOATING
C610 A2c 0 1.6834f **FLOATING
C611 xor_2 0 1.63601f **FLOATING
C612 DEC_D0_NAND 0 0.511796f **FLOATING
C613 ander_node_5 0 0.248064f **FLOATING
C614 ander_node_6 0 0.248064f **FLOATING
C615 ander_node_7 0 0.248064f **FLOATING
C616 S1c 0 4.36861f **FLOATING
C617 S0c 0 5.09312f **FLOATING
C618 ander_node_8 0 0.248064f **FLOATING
C619 and_b0e_nand 0 0.52029f **FLOATING
C620 and_b1e_nand 0 0.52029f **FLOATING
C621 and_b2e_nand 0 0.52029f **FLOATING
C622 and_b3e_nand 0 0.52029f **FLOATING
C623 B0 0 27.8381f **FLOATING
C624 B1 0 23.611198f **FLOATING
C625 B2 0 18.705599f **FLOATING
C626 B3 0 11.262401f **FLOATING
C627 ander_node_12 0 0.248064f **FLOATING
C628 ander_node_11 0 0.248064f **FLOATING
C629 ander_node_10 0 0.248064f **FLOATING
C630 ander_node_9 0 0.248064f **FLOATING
C631 A0_and_B0 0 0.075352f **FLOATING
C632 A1_and_B1 0 0.075352f **FLOATING
C633 A2_and_B2 0 0.075352f **FLOATING
C634 A3_and_B3 0 0.075352f **FLOATING
C635 ander_node_4 0 0.248064f **FLOATING
C636 ander_node_3 0 0.248064f **FLOATING
C637 ander_node_2 0 0.248064f **FLOATING
C638 ander_node_1 0 0.248064f **FLOATING
C639 A0_and_B0_nand 0 0.52029f **FLOATING
C640 A1_and_B1_nand 0 0.52029f **FLOATING
C641 A2_and_B2_nand 0 0.52029f **FLOATING
C642 A3_and_B3_nand 0 0.52029f **FLOATING
C643 and_b0e 0 3.10166f **FLOATING
C644 and_a0e 0 3.54193f **FLOATING
C645 and_b1e 0 3.64923f **FLOATING
C646 and_a1e 0 5.29932f **FLOATING
C647 and_b2e 0 3.87059f **FLOATING
C648 and_a2e 0 5.463779f **FLOATING
C649 and_b3e 0 3.78326f **FLOATING
C650 and_a3e 0 9.534531f **FLOATING
C651 and_a0e_nand 0 0.52029f **FLOATING
C652 and_a1e_nand 0 0.52029f **FLOATING
C653 and_a2e_nand 0 0.52029f **FLOATING
C654 and_a3e_nand 0 0.52029f **FLOATING
C655 A_greater_B_node_1 0 0.248064f **FLOATING
C656 compare_B3e 0 16.0881f **FLOATING
C657 A0 0 24.168f **FLOATING
C658 A1 0 20.3698f **FLOATING
C659 A2 0 13.563f **FLOATING
C660 D3 0 23.219599f **FLOATING
C661 A3 0 11.0655f **FLOATING
C662 A3_nand_B3c 0 0.52029f **FLOATING
C663 compare_A2e 0 14.2568f **FLOATING
C664 A3c 0 1.6834f **FLOATING
C665 compare_A3e 0 12.8447f **FLOATING
C666 xor_1 0 1.64089f **FLOATING
C667 B3c 0 12.7175f **FLOATING
C668 A3_eq_B3_A2_gt_B2_c 0 0.59518f **FLOATING
C669 compare_A1e 0 15.1418f **FLOATING
C670 a_754_699# 0 0.388565f **FLOATING
C671 A3_eq_B3_A2_eq_B2_A1_gt_B1_c 0 0.617397f **FLOATING
C672 B2c 0 7.22845f **FLOATING
C673 B1c 0 7.55881f **FLOATING
C674 A3e_xnor_B3e 0 19.5984f **FLOATING
C675 a_706_699# 0 0.388565f **FLOATING
C676 a_690_700# 0 0.38028f **FLOATING
C677 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c 0 0.644677f **FLOATING
C678 A2e_xnor_B2e 0 9.465691f **FLOATING
C679 A3_and_B3c 0 3.03158f **FLOATING
C680 A3_eq_B3_A2_gt_B2 0 2.92765f **FLOATING
C681 A3_eq_B3_A2_eq_B2_A1_gt_B1 0 1.909f **FLOATING
C682 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0 0 2.4789f **FLOATING
C683 A_GT_B 0 0.421262f **FLOATING
C684 A_GT_B_c 0 0.668379f **FLOATING
C685 gnd 0 68.3142f **FLOATING
C686 A_LS_B_node_1 0 0.248064f **FLOATING
C687 A_LS_B 0 0.101396f **FLOATING
C688 A_LS_B_nand 0 0.52029f **FLOATING
C689 a_840_939# 0 1.40121f **FLOATING
C690 A_equal_B_c 0 18.6104f **FLOATING
C691 vdd 0 0.153228p **FLOATING
