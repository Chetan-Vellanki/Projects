magic
tech scmos
timestamp 1701523321
<< nwell >>
rect 863 1568 909 1587
rect 923 1584 984 1601
rect 647 1505 731 1506
rect 647 1486 798 1505
rect 809 1487 855 1506
rect 647 1476 752 1486
rect 666 1302 776 1303
rect 855 1302 954 1303
rect 620 1283 776 1302
rect 809 1283 954 1302
rect 967 1283 1013 1302
rect 674 1274 776 1283
rect 855 1274 954 1283
rect 1020 1270 1097 1302
rect 297 1266 361 1267
rect 186 1247 232 1266
rect 257 1247 361 1266
rect 1125 1265 1171 1284
rect 1185 1281 1246 1298
rect 308 1240 361 1247
rect 309 1239 361 1240
rect 376 1200 443 1228
rect 458 1204 504 1223
rect 294 1044 358 1045
rect 183 1025 229 1044
rect 254 1025 358 1044
rect 305 1018 358 1025
rect 678 1019 724 1038
rect 738 1035 799 1052
rect 825 1019 871 1038
rect 885 1035 946 1052
rect 306 1017 358 1018
rect 971 1017 1017 1036
rect 1031 1033 1092 1050
rect 1107 1017 1153 1036
rect 1167 1033 1228 1050
rect 380 1006 403 1011
rect 373 978 440 1006
rect 455 982 501 1001
rect 669 912 715 931
rect 729 928 790 945
rect 814 911 860 930
rect 874 927 935 944
rect 963 909 1009 928
rect 1023 925 1084 942
rect 1107 909 1153 928
rect 1167 925 1228 942
rect 49 871 147 872
rect 3 852 147 871
rect 297 859 361 860
rect 49 843 147 852
rect 161 840 232 859
rect 257 840 361 859
rect 308 833 361 840
rect 309 832 361 833
rect 388 824 406 826
rect 383 821 406 824
rect 376 793 443 821
rect 458 797 504 816
rect 297 684 361 685
rect 186 665 232 684
rect 257 665 361 684
rect 308 658 361 665
rect 309 657 361 658
rect 379 646 406 651
rect 376 618 443 646
rect 458 622 504 641
<< ntransistor >>
rect 936 1561 941 1566
rect 959 1561 964 1566
rect 878 1553 883 1558
rect 778 1471 783 1476
rect 835 1472 840 1477
rect 669 1453 674 1458
rect 685 1453 690 1458
rect 701 1453 706 1458
rect 717 1453 722 1458
rect 635 1268 640 1273
rect 824 1268 829 1273
rect 982 1268 987 1273
rect 406 1250 411 1255
rect 424 1250 429 1255
rect 690 1252 695 1257
rect 706 1252 711 1257
rect 722 1252 727 1257
rect 738 1252 743 1257
rect 754 1252 759 1257
rect 883 1252 888 1257
rect 899 1252 904 1257
rect 915 1252 920 1257
rect 931 1252 936 1257
rect 212 1232 217 1237
rect 272 1232 277 1237
rect 1045 1251 1050 1256
rect 1061 1251 1066 1256
rect 1077 1251 1082 1256
rect 1198 1258 1203 1263
rect 1221 1258 1226 1263
rect 1140 1250 1145 1255
rect 323 1211 328 1216
rect 341 1211 346 1216
rect 484 1189 489 1194
rect 403 1028 408 1033
rect 421 1028 426 1033
rect 209 1010 214 1015
rect 269 1010 274 1015
rect 320 989 325 994
rect 338 989 343 994
rect 751 1012 756 1017
rect 774 1012 779 1017
rect 693 1004 698 1009
rect 898 1012 903 1017
rect 921 1012 926 1017
rect 840 1004 845 1009
rect 1044 1010 1049 1015
rect 1067 1010 1072 1015
rect 986 1002 991 1007
rect 1180 1010 1185 1015
rect 1203 1010 1208 1015
rect 1122 1002 1127 1007
rect 481 967 486 972
rect 742 905 747 910
rect 765 905 770 910
rect 684 897 689 902
rect 887 904 892 909
rect 910 904 915 909
rect 829 896 834 901
rect 1036 902 1041 907
rect 1059 902 1064 907
rect 978 894 983 899
rect 1180 902 1185 907
rect 1203 902 1208 907
rect 1122 894 1127 899
rect 18 837 23 842
rect 406 843 411 848
rect 424 843 429 848
rect 77 821 82 826
rect 93 821 98 826
rect 109 821 114 826
rect 125 821 130 826
rect 212 825 217 830
rect 272 825 277 830
rect 323 804 328 809
rect 341 804 346 809
rect 484 782 489 787
rect 406 668 411 673
rect 424 668 429 673
rect 212 650 217 655
rect 272 650 277 655
rect 323 629 328 634
rect 341 629 346 634
rect 484 607 489 612
<< ptransistor >>
rect 936 1590 941 1595
rect 959 1590 964 1595
rect 878 1575 883 1580
rect 669 1489 674 1494
rect 685 1489 690 1494
rect 701 1489 706 1494
rect 717 1489 722 1494
rect 778 1493 783 1498
rect 835 1494 840 1499
rect 635 1290 640 1295
rect 690 1286 695 1291
rect 706 1286 711 1291
rect 722 1286 727 1291
rect 738 1286 743 1291
rect 754 1286 759 1291
rect 824 1290 829 1295
rect 212 1254 217 1259
rect 272 1254 277 1259
rect 883 1286 888 1291
rect 899 1286 904 1291
rect 915 1286 920 1291
rect 931 1286 936 1291
rect 982 1290 987 1295
rect 1045 1285 1050 1290
rect 1061 1285 1066 1290
rect 1077 1285 1082 1290
rect 1198 1287 1203 1292
rect 1221 1287 1226 1292
rect 323 1250 328 1255
rect 341 1250 346 1255
rect 1140 1272 1145 1277
rect 406 1211 411 1216
rect 424 1211 429 1216
rect 484 1211 489 1216
rect 209 1032 214 1037
rect 269 1032 274 1037
rect 751 1041 756 1046
rect 774 1041 779 1046
rect 898 1041 903 1046
rect 921 1041 926 1046
rect 320 1028 325 1033
rect 338 1028 343 1033
rect 693 1026 698 1031
rect 840 1026 845 1031
rect 1044 1039 1049 1044
rect 1067 1039 1072 1044
rect 1180 1039 1185 1044
rect 1203 1039 1208 1044
rect 986 1024 991 1029
rect 403 989 408 994
rect 421 989 426 994
rect 481 989 486 994
rect 1122 1024 1127 1029
rect 742 934 747 939
rect 765 934 770 939
rect 684 919 689 924
rect 887 933 892 938
rect 910 933 915 938
rect 829 918 834 923
rect 1036 931 1041 936
rect 1059 931 1064 936
rect 1180 931 1185 936
rect 1203 931 1208 936
rect 978 916 983 921
rect 1122 916 1127 921
rect 18 859 23 864
rect 77 855 82 860
rect 93 855 98 860
rect 109 855 114 860
rect 125 855 130 860
rect 212 847 217 852
rect 272 847 277 852
rect 323 843 328 848
rect 341 843 346 848
rect 406 804 411 809
rect 424 804 429 809
rect 484 804 489 809
rect 212 672 217 677
rect 272 672 277 677
rect 323 668 328 673
rect 341 668 346 673
rect 406 629 411 634
rect 424 629 429 634
rect 484 629 489 634
<< ndiffusion >>
rect 934 1561 936 1566
rect 941 1561 943 1566
rect 957 1561 959 1566
rect 964 1561 966 1566
rect 875 1553 878 1558
rect 883 1553 885 1558
rect 776 1471 778 1476
rect 783 1471 786 1476
rect 833 1472 835 1477
rect 840 1472 843 1477
rect 666 1453 669 1458
rect 674 1453 677 1458
rect 682 1453 685 1458
rect 690 1453 693 1458
rect 698 1453 701 1458
rect 706 1453 709 1458
rect 714 1453 717 1458
rect 722 1453 725 1458
rect 632 1268 635 1273
rect 640 1268 642 1273
rect 821 1268 824 1273
rect 829 1268 831 1273
rect 979 1268 982 1273
rect 987 1268 989 1273
rect 403 1250 406 1255
rect 411 1250 424 1255
rect 429 1250 432 1255
rect 687 1252 690 1257
rect 695 1252 706 1257
rect 711 1252 722 1257
rect 727 1252 738 1257
rect 743 1252 754 1257
rect 759 1252 762 1257
rect 881 1252 883 1257
rect 888 1252 899 1257
rect 904 1252 915 1257
rect 920 1252 931 1257
rect 936 1252 939 1257
rect 210 1232 212 1237
rect 217 1232 220 1237
rect 269 1232 272 1237
rect 277 1232 279 1237
rect 1039 1251 1045 1256
rect 1050 1251 1061 1256
rect 1066 1251 1077 1256
rect 1082 1251 1085 1256
rect 1196 1258 1198 1263
rect 1203 1258 1205 1263
rect 1219 1258 1221 1263
rect 1226 1258 1228 1263
rect 1137 1250 1140 1255
rect 1145 1250 1147 1255
rect 320 1211 323 1216
rect 328 1211 341 1216
rect 346 1211 349 1216
rect 482 1189 484 1194
rect 489 1189 492 1194
rect 400 1028 403 1033
rect 408 1028 421 1033
rect 426 1028 429 1033
rect 207 1010 209 1015
rect 214 1010 217 1015
rect 266 1010 269 1015
rect 274 1010 276 1015
rect 317 989 320 994
rect 325 989 338 994
rect 343 989 346 994
rect 749 1012 751 1017
rect 756 1012 758 1017
rect 772 1012 774 1017
rect 779 1012 781 1017
rect 690 1004 693 1009
rect 698 1004 700 1009
rect 896 1012 898 1017
rect 903 1012 905 1017
rect 919 1012 921 1017
rect 926 1012 928 1017
rect 837 1004 840 1009
rect 845 1004 847 1009
rect 1042 1010 1044 1015
rect 1049 1010 1051 1015
rect 1065 1010 1067 1015
rect 1072 1010 1074 1015
rect 983 1002 986 1007
rect 991 1002 993 1007
rect 1178 1010 1180 1015
rect 1185 1010 1187 1015
rect 1201 1010 1203 1015
rect 1208 1010 1210 1015
rect 1119 1002 1122 1007
rect 1127 1002 1129 1007
rect 479 967 481 972
rect 486 967 489 972
rect 740 905 742 910
rect 747 905 749 910
rect 763 905 765 910
rect 770 905 772 910
rect 681 897 684 902
rect 689 897 691 902
rect 885 904 887 909
rect 892 904 894 909
rect 908 904 910 909
rect 915 904 917 909
rect 826 896 829 901
rect 834 896 836 901
rect 1034 902 1036 907
rect 1041 902 1043 907
rect 1057 902 1059 907
rect 1064 902 1066 907
rect 975 894 978 899
rect 983 894 985 899
rect 1178 902 1180 907
rect 1185 902 1187 907
rect 1201 902 1203 907
rect 1208 902 1210 907
rect 1119 894 1122 899
rect 1127 894 1129 899
rect 15 837 18 842
rect 23 837 25 842
rect 403 843 406 848
rect 411 843 424 848
rect 429 843 432 848
rect 75 821 77 826
rect 82 821 93 826
rect 98 821 109 826
rect 114 821 125 826
rect 130 821 133 826
rect 210 825 212 830
rect 217 825 220 830
rect 269 825 272 830
rect 277 825 279 830
rect 320 804 323 809
rect 328 804 341 809
rect 346 804 349 809
rect 482 782 484 787
rect 489 782 492 787
rect 403 668 406 673
rect 411 668 424 673
rect 429 668 432 673
rect 210 650 212 655
rect 217 650 220 655
rect 269 650 272 655
rect 277 650 279 655
rect 320 629 323 634
rect 328 629 341 634
rect 346 629 349 634
rect 482 607 484 612
rect 489 607 492 612
<< pdiffusion >>
rect 934 1590 936 1595
rect 941 1590 947 1595
rect 952 1590 959 1595
rect 964 1590 966 1595
rect 875 1575 878 1580
rect 883 1575 885 1580
rect 666 1489 669 1494
rect 674 1489 685 1494
rect 690 1489 701 1494
rect 706 1489 717 1494
rect 722 1489 725 1494
rect 776 1493 778 1498
rect 783 1493 786 1498
rect 833 1494 835 1499
rect 840 1494 843 1499
rect 632 1290 635 1295
rect 640 1290 642 1295
rect 687 1286 690 1291
rect 695 1286 698 1291
rect 703 1286 706 1291
rect 711 1286 714 1291
rect 719 1286 722 1291
rect 727 1286 730 1291
rect 735 1286 738 1291
rect 743 1286 746 1291
rect 751 1286 754 1291
rect 759 1286 762 1291
rect 821 1290 824 1295
rect 829 1290 831 1295
rect 210 1254 212 1259
rect 217 1254 220 1259
rect 269 1254 272 1259
rect 277 1254 279 1259
rect 880 1286 883 1291
rect 888 1286 891 1291
rect 896 1286 899 1291
rect 904 1286 907 1291
rect 912 1286 915 1291
rect 920 1286 923 1291
rect 928 1286 931 1291
rect 936 1286 939 1291
rect 979 1290 982 1295
rect 987 1290 989 1295
rect 1042 1285 1045 1290
rect 1050 1285 1053 1290
rect 1058 1285 1061 1290
rect 1066 1285 1069 1290
rect 1074 1285 1077 1290
rect 1082 1285 1085 1290
rect 1196 1287 1198 1292
rect 1203 1287 1209 1292
rect 1214 1287 1221 1292
rect 1226 1287 1228 1292
rect 320 1250 323 1255
rect 328 1250 341 1255
rect 346 1250 349 1255
rect 1137 1272 1140 1277
rect 1145 1272 1147 1277
rect 403 1211 406 1216
rect 411 1211 424 1216
rect 429 1211 432 1216
rect 482 1211 484 1216
rect 489 1211 492 1216
rect 207 1032 209 1037
rect 214 1032 217 1037
rect 266 1032 269 1037
rect 274 1032 276 1037
rect 749 1041 751 1046
rect 756 1041 762 1046
rect 767 1041 774 1046
rect 779 1041 781 1046
rect 896 1041 898 1046
rect 903 1041 909 1046
rect 914 1041 921 1046
rect 926 1041 928 1046
rect 317 1028 320 1033
rect 325 1028 338 1033
rect 343 1028 346 1033
rect 690 1026 693 1031
rect 698 1026 700 1031
rect 837 1026 840 1031
rect 845 1026 847 1031
rect 1042 1039 1044 1044
rect 1049 1039 1055 1044
rect 1060 1039 1067 1044
rect 1072 1039 1074 1044
rect 1178 1039 1180 1044
rect 1185 1039 1191 1044
rect 1196 1039 1203 1044
rect 1208 1039 1210 1044
rect 983 1024 986 1029
rect 991 1024 993 1029
rect 400 989 403 994
rect 408 989 421 994
rect 426 989 429 994
rect 479 989 481 994
rect 486 989 489 994
rect 1119 1024 1122 1029
rect 1127 1024 1129 1029
rect 740 934 742 939
rect 747 934 753 939
rect 758 934 765 939
rect 770 934 772 939
rect 681 919 684 924
rect 689 919 691 924
rect 885 933 887 938
rect 892 933 898 938
rect 903 933 910 938
rect 915 933 917 938
rect 826 918 829 923
rect 834 918 836 923
rect 1034 931 1036 936
rect 1041 931 1047 936
rect 1052 931 1059 936
rect 1064 931 1066 936
rect 1178 931 1180 936
rect 1185 931 1191 936
rect 1196 931 1203 936
rect 1208 931 1210 936
rect 975 916 978 921
rect 983 916 985 921
rect 1119 916 1122 921
rect 1127 916 1129 921
rect 15 859 18 864
rect 23 859 25 864
rect 74 855 77 860
rect 82 855 85 860
rect 90 855 93 860
rect 98 855 101 860
rect 106 855 109 860
rect 114 855 117 860
rect 122 855 125 860
rect 130 855 133 860
rect 210 847 212 852
rect 217 847 220 852
rect 269 847 272 852
rect 277 847 279 852
rect 320 843 323 848
rect 328 843 341 848
rect 346 843 349 848
rect 403 804 406 809
rect 411 804 424 809
rect 429 804 432 809
rect 482 804 484 809
rect 489 804 492 809
rect 210 672 212 677
rect 217 672 220 677
rect 269 672 272 677
rect 277 672 279 677
rect 320 668 323 673
rect 328 668 341 673
rect 346 668 349 673
rect 403 629 406 634
rect 411 629 424 634
rect 429 629 432 634
rect 482 629 484 634
rect 489 629 492 634
<< ndcontact >>
rect 929 1561 934 1566
rect 943 1561 947 1566
rect 953 1561 957 1566
rect 966 1561 971 1566
rect 870 1553 875 1558
rect 885 1553 890 1558
rect 771 1471 776 1476
rect 786 1471 791 1476
rect 828 1472 833 1477
rect 843 1472 848 1477
rect 661 1453 666 1458
rect 677 1453 682 1458
rect 693 1453 698 1458
rect 709 1453 714 1458
rect 725 1453 730 1458
rect 627 1268 632 1273
rect 642 1268 647 1273
rect 816 1268 821 1273
rect 831 1268 836 1273
rect 974 1268 979 1273
rect 989 1268 994 1273
rect 398 1250 403 1255
rect 432 1250 437 1255
rect 682 1252 687 1257
rect 762 1252 767 1257
rect 876 1252 881 1257
rect 939 1252 944 1257
rect 205 1232 210 1237
rect 220 1232 225 1237
rect 264 1232 269 1237
rect 279 1232 284 1237
rect 1034 1251 1039 1256
rect 1085 1251 1090 1256
rect 1191 1258 1196 1263
rect 1205 1258 1209 1263
rect 1215 1258 1219 1263
rect 1228 1258 1233 1263
rect 1132 1250 1137 1255
rect 1147 1250 1152 1255
rect 315 1211 320 1216
rect 349 1211 354 1216
rect 477 1189 482 1194
rect 492 1189 497 1194
rect 395 1028 400 1033
rect 429 1028 434 1033
rect 202 1010 207 1015
rect 217 1010 222 1015
rect 261 1010 266 1015
rect 276 1010 281 1015
rect 312 989 317 994
rect 346 989 351 994
rect 744 1012 749 1017
rect 758 1012 762 1017
rect 768 1012 772 1017
rect 781 1012 786 1017
rect 685 1004 690 1009
rect 700 1004 705 1009
rect 891 1012 896 1017
rect 905 1012 909 1017
rect 915 1012 919 1017
rect 928 1012 933 1017
rect 832 1004 837 1009
rect 847 1004 852 1009
rect 1037 1010 1042 1015
rect 1051 1010 1055 1015
rect 1061 1010 1065 1015
rect 1074 1010 1079 1015
rect 978 1002 983 1007
rect 993 1002 998 1007
rect 1173 1010 1178 1015
rect 1187 1010 1191 1015
rect 1197 1010 1201 1015
rect 1210 1010 1215 1015
rect 1114 1002 1119 1007
rect 1129 1002 1134 1007
rect 474 967 479 972
rect 489 967 494 972
rect 735 905 740 910
rect 749 905 753 910
rect 759 905 763 910
rect 772 905 777 910
rect 676 897 681 902
rect 691 897 696 902
rect 880 904 885 909
rect 894 904 898 909
rect 904 904 908 909
rect 917 904 922 909
rect 821 896 826 901
rect 836 896 841 901
rect 1029 902 1034 907
rect 1043 902 1047 907
rect 1053 902 1057 907
rect 1066 902 1071 907
rect 970 894 975 899
rect 985 894 990 899
rect 1173 902 1178 907
rect 1187 902 1191 907
rect 1197 902 1201 907
rect 1210 902 1215 907
rect 1114 894 1119 899
rect 1129 894 1134 899
rect 10 837 15 842
rect 25 837 30 842
rect 398 843 403 848
rect 432 843 437 848
rect 70 821 75 826
rect 133 821 138 826
rect 205 825 210 830
rect 220 825 225 830
rect 264 825 269 830
rect 279 825 284 830
rect 315 804 320 809
rect 349 804 354 809
rect 477 782 482 787
rect 492 782 497 787
rect 398 668 403 673
rect 432 668 437 673
rect 205 650 210 655
rect 220 650 225 655
rect 264 650 269 655
rect 279 650 284 655
rect 315 629 320 634
rect 349 629 354 634
rect 477 607 482 612
rect 492 607 497 612
<< pdcontact >>
rect 929 1590 934 1595
rect 947 1590 952 1595
rect 966 1590 971 1595
rect 870 1575 875 1580
rect 885 1575 890 1580
rect 661 1489 666 1494
rect 725 1489 730 1494
rect 771 1493 776 1498
rect 786 1493 791 1498
rect 828 1494 833 1499
rect 843 1494 848 1499
rect 627 1290 632 1295
rect 642 1290 647 1295
rect 682 1286 687 1291
rect 698 1286 703 1291
rect 714 1286 719 1291
rect 730 1286 735 1291
rect 746 1286 751 1291
rect 762 1286 767 1291
rect 816 1290 821 1295
rect 831 1290 836 1295
rect 205 1254 210 1259
rect 220 1254 225 1259
rect 264 1254 269 1259
rect 279 1254 284 1259
rect 875 1286 880 1291
rect 891 1286 896 1291
rect 907 1286 912 1291
rect 923 1286 928 1291
rect 939 1286 944 1291
rect 974 1290 979 1295
rect 989 1290 994 1295
rect 1037 1285 1042 1290
rect 1053 1285 1058 1290
rect 1069 1285 1074 1290
rect 1085 1285 1090 1290
rect 1191 1287 1196 1292
rect 1209 1287 1214 1292
rect 1228 1287 1233 1292
rect 315 1250 320 1255
rect 349 1250 354 1255
rect 1132 1272 1137 1277
rect 1147 1272 1152 1277
rect 398 1211 403 1216
rect 432 1211 437 1216
rect 477 1211 482 1216
rect 492 1211 497 1216
rect 202 1032 207 1037
rect 217 1032 222 1037
rect 261 1032 266 1037
rect 276 1032 281 1037
rect 744 1041 749 1046
rect 762 1041 767 1046
rect 781 1041 786 1046
rect 891 1041 896 1046
rect 909 1041 914 1046
rect 928 1041 933 1046
rect 312 1028 317 1033
rect 346 1028 351 1033
rect 685 1026 690 1031
rect 700 1026 705 1031
rect 832 1026 837 1031
rect 847 1026 852 1031
rect 1037 1039 1042 1044
rect 1055 1039 1060 1044
rect 1074 1039 1079 1044
rect 1173 1039 1178 1044
rect 1191 1039 1196 1044
rect 1210 1039 1215 1044
rect 978 1024 983 1029
rect 993 1024 998 1029
rect 395 989 400 994
rect 429 989 434 994
rect 474 989 479 994
rect 489 989 494 994
rect 1114 1024 1119 1029
rect 1129 1024 1134 1029
rect 735 934 740 939
rect 753 934 758 939
rect 772 934 777 939
rect 676 919 681 924
rect 691 919 696 924
rect 880 933 885 938
rect 898 933 903 938
rect 917 933 922 938
rect 821 918 826 923
rect 836 918 841 923
rect 1029 931 1034 936
rect 1047 931 1052 936
rect 1066 931 1071 936
rect 1173 931 1178 936
rect 1191 931 1196 936
rect 1210 931 1215 936
rect 970 916 975 921
rect 985 916 990 921
rect 1114 916 1119 921
rect 1129 916 1134 921
rect 10 859 15 864
rect 25 859 30 864
rect 69 855 74 860
rect 85 855 90 860
rect 101 855 106 860
rect 117 855 122 860
rect 133 855 138 860
rect 205 847 210 852
rect 220 847 225 852
rect 264 847 269 852
rect 279 847 284 852
rect 315 843 320 848
rect 349 843 354 848
rect 398 804 403 809
rect 432 804 437 809
rect 477 804 482 809
rect 492 804 497 809
rect 205 672 210 677
rect 220 672 225 677
rect 264 672 269 677
rect 279 672 284 677
rect 315 668 320 673
rect 349 668 354 673
rect 398 629 403 634
rect 432 629 437 634
rect 477 629 482 634
rect 492 629 497 634
<< nsubstratencontact >>
rect 975 1590 980 1595
rect 897 1575 902 1580
rect 737 1489 742 1494
rect 759 1493 764 1498
rect 816 1494 821 1499
rect 654 1290 659 1295
rect 843 1290 848 1295
rect 193 1254 198 1259
rect 291 1254 296 1259
rect 863 1286 868 1291
rect 1001 1290 1006 1295
rect 1027 1285 1032 1290
rect 1237 1287 1242 1292
rect 303 1250 308 1255
rect 1159 1272 1164 1277
rect 383 1209 389 1215
rect 465 1211 470 1216
rect 190 1032 195 1037
rect 288 1032 293 1037
rect 790 1041 795 1046
rect 937 1041 942 1046
rect 300 1028 305 1033
rect 712 1026 717 1031
rect 859 1026 864 1031
rect 1083 1039 1088 1044
rect 1219 1039 1224 1044
rect 1005 1024 1010 1029
rect 380 990 386 995
rect 462 989 467 994
rect 1141 1024 1146 1029
rect 781 934 786 939
rect 703 919 708 924
rect 926 933 931 938
rect 848 918 853 923
rect 1075 931 1080 936
rect 1219 931 1224 936
rect 997 916 1002 921
rect 1141 916 1146 921
rect 37 859 42 864
rect 57 855 62 860
rect 168 847 173 852
rect 291 847 296 852
rect 303 843 308 848
rect 383 802 388 808
rect 465 804 470 809
rect 193 672 198 677
rect 291 672 296 677
rect 303 668 308 673
rect 383 629 388 634
rect 465 629 470 634
<< polysilicon >>
rect 936 1595 941 1609
rect 959 1595 964 1609
rect 878 1580 883 1583
rect 878 1566 883 1575
rect 936 1566 941 1590
rect 959 1566 964 1590
rect 878 1562 882 1566
rect 878 1558 883 1562
rect 878 1548 883 1553
rect 936 1542 941 1561
rect 959 1542 964 1561
rect 778 1498 783 1501
rect 835 1499 840 1502
rect 669 1494 674 1497
rect 685 1494 690 1497
rect 701 1494 706 1497
rect 717 1494 722 1497
rect 669 1458 674 1489
rect 685 1458 690 1489
rect 701 1458 706 1489
rect 717 1458 722 1489
rect 778 1484 783 1493
rect 835 1485 840 1494
rect 779 1480 783 1484
rect 836 1481 840 1485
rect 778 1476 783 1480
rect 835 1477 840 1481
rect 778 1466 783 1471
rect 835 1467 840 1472
rect 669 1442 674 1453
rect 685 1442 690 1453
rect 701 1442 706 1453
rect 717 1443 722 1453
rect 635 1295 640 1298
rect 690 1291 695 1295
rect 706 1291 711 1295
rect 722 1291 727 1310
rect 738 1291 743 1310
rect 824 1295 829 1298
rect 754 1291 759 1295
rect 635 1281 640 1290
rect 883 1291 888 1310
rect 899 1291 904 1310
rect 915 1291 920 1295
rect 931 1291 936 1310
rect 982 1295 987 1298
rect 341 1276 379 1277
rect 635 1277 639 1281
rect 384 1276 429 1277
rect 341 1272 429 1276
rect 635 1273 640 1277
rect 212 1259 217 1262
rect 272 1259 277 1262
rect 323 1255 328 1259
rect 341 1255 346 1272
rect 406 1255 411 1259
rect 424 1255 429 1272
rect 635 1263 640 1268
rect 690 1257 695 1286
rect 706 1257 711 1286
rect 722 1257 727 1286
rect 738 1257 743 1286
rect 754 1257 759 1286
rect 824 1281 829 1290
rect 1045 1290 1050 1295
rect 1061 1290 1066 1312
rect 1077 1290 1082 1310
rect 1198 1292 1203 1306
rect 1221 1292 1226 1306
rect 824 1277 828 1281
rect 824 1273 829 1277
rect 824 1263 829 1268
rect 883 1257 888 1286
rect 899 1257 904 1286
rect 915 1257 920 1286
rect 931 1257 936 1286
rect 982 1281 987 1290
rect 982 1277 986 1281
rect 982 1273 987 1277
rect 982 1263 987 1268
rect 212 1245 217 1254
rect 213 1241 217 1245
rect 212 1237 217 1241
rect 272 1245 277 1254
rect 1045 1256 1050 1285
rect 1061 1256 1066 1285
rect 1077 1256 1082 1285
rect 1140 1277 1145 1280
rect 1140 1263 1145 1272
rect 1198 1263 1203 1287
rect 1221 1263 1226 1287
rect 1140 1259 1144 1263
rect 272 1241 276 1245
rect 272 1237 277 1241
rect 323 1238 328 1250
rect 341 1246 346 1250
rect 406 1238 411 1250
rect 424 1246 429 1250
rect 324 1233 346 1238
rect 406 1233 429 1238
rect 690 1233 695 1252
rect 212 1227 217 1232
rect 272 1227 277 1232
rect 304 1221 328 1226
rect 304 1213 309 1221
rect 323 1216 328 1221
rect 341 1216 346 1233
rect 406 1216 411 1220
rect 424 1216 429 1233
rect 706 1232 711 1252
rect 722 1235 727 1252
rect 738 1235 743 1252
rect 754 1232 759 1252
rect 883 1245 888 1252
rect 899 1245 904 1252
rect 915 1235 920 1252
rect 931 1235 936 1252
rect 1140 1255 1145 1259
rect 1045 1236 1050 1251
rect 1061 1237 1066 1251
rect 1077 1237 1082 1251
rect 1140 1245 1145 1250
rect 1198 1239 1203 1258
rect 1221 1239 1226 1258
rect 484 1216 489 1219
rect 323 1193 328 1211
rect 341 1205 346 1211
rect 406 1193 411 1211
rect 323 1188 411 1193
rect 424 1176 429 1211
rect 484 1202 489 1211
rect 485 1198 489 1202
rect 484 1194 489 1198
rect 484 1184 489 1189
rect 338 1054 376 1055
rect 381 1054 426 1055
rect 338 1050 426 1054
rect 209 1037 214 1040
rect 269 1037 274 1040
rect 320 1033 325 1037
rect 338 1033 343 1050
rect 403 1033 408 1037
rect 421 1033 426 1050
rect 751 1046 756 1060
rect 774 1046 779 1060
rect 898 1046 903 1060
rect 921 1046 926 1060
rect 1044 1044 1049 1058
rect 1067 1044 1072 1058
rect 1180 1044 1185 1058
rect 1203 1044 1208 1058
rect 209 1023 214 1032
rect 210 1019 214 1023
rect 209 1015 214 1019
rect 269 1023 274 1032
rect 693 1031 698 1034
rect 269 1019 273 1023
rect 269 1015 274 1019
rect 320 1016 325 1028
rect 338 1024 343 1028
rect 403 1016 408 1028
rect 421 1024 426 1028
rect 693 1017 698 1026
rect 751 1017 756 1041
rect 774 1017 779 1041
rect 840 1031 845 1034
rect 840 1017 845 1026
rect 898 1017 903 1041
rect 921 1017 926 1041
rect 986 1029 991 1032
rect 321 1011 343 1016
rect 403 1011 426 1016
rect 209 1005 214 1010
rect 269 1005 274 1010
rect 301 999 325 1004
rect 301 991 306 999
rect 320 994 325 999
rect 338 994 343 1011
rect 403 994 408 998
rect 421 994 426 1011
rect 693 1013 697 1017
rect 693 1009 698 1013
rect 840 1013 844 1017
rect 693 999 698 1004
rect 481 994 486 997
rect 751 993 756 1012
rect 320 971 325 989
rect 338 983 343 989
rect 403 971 408 989
rect 320 966 408 971
rect 421 954 426 989
rect 481 980 486 989
rect 774 993 779 1012
rect 840 1009 845 1013
rect 986 1015 991 1024
rect 1044 1015 1049 1039
rect 1067 1015 1072 1039
rect 1122 1029 1127 1032
rect 1122 1015 1127 1024
rect 1180 1015 1185 1039
rect 1203 1015 1208 1039
rect 840 999 845 1004
rect 898 993 903 1012
rect 921 993 926 1012
rect 986 1011 990 1015
rect 986 1007 991 1011
rect 1122 1011 1126 1015
rect 986 997 991 1002
rect 1044 991 1049 1010
rect 1067 991 1072 1010
rect 1122 1007 1127 1011
rect 1122 997 1127 1002
rect 1180 991 1185 1010
rect 1203 991 1208 1010
rect 482 976 486 980
rect 481 972 486 976
rect 481 962 486 967
rect 742 939 747 953
rect 765 939 770 953
rect 887 938 892 952
rect 910 938 915 952
rect 684 924 689 927
rect 684 910 689 919
rect 742 910 747 934
rect 765 910 770 934
rect 1036 936 1041 950
rect 1059 936 1064 950
rect 1180 936 1185 950
rect 1203 936 1208 950
rect 829 923 834 926
rect 684 906 688 910
rect 684 902 689 906
rect 829 909 834 918
rect 887 909 892 933
rect 910 909 915 933
rect 978 921 983 924
rect 829 905 833 909
rect 684 892 689 897
rect 742 886 747 905
rect 765 886 770 905
rect 829 901 834 905
rect 978 907 983 916
rect 1036 907 1041 931
rect 1059 907 1064 931
rect 1122 921 1127 924
rect 1122 907 1127 916
rect 1180 907 1185 931
rect 1203 907 1208 931
rect 829 891 834 896
rect 887 885 892 904
rect 910 885 915 904
rect 978 903 982 907
rect 978 899 983 903
rect 1122 903 1126 907
rect 978 889 983 894
rect 1036 883 1041 902
rect 18 864 23 867
rect 77 860 82 879
rect 93 860 98 879
rect 1059 883 1064 902
rect 1122 899 1127 903
rect 1122 889 1127 894
rect 1180 883 1185 902
rect 1203 883 1208 902
rect 341 869 379 870
rect 384 869 429 870
rect 341 865 429 869
rect 109 860 114 864
rect 125 860 130 864
rect 18 850 23 859
rect 18 846 22 850
rect 18 842 23 846
rect 18 832 23 837
rect 77 826 82 855
rect 93 826 98 855
rect 109 826 114 855
rect 125 826 130 855
rect 212 852 217 855
rect 272 852 277 855
rect 323 848 328 852
rect 341 848 346 865
rect 406 848 411 852
rect 424 848 429 865
rect 212 838 217 847
rect 213 834 217 838
rect 212 830 217 834
rect 272 838 277 847
rect 272 834 276 838
rect 272 830 277 834
rect 323 831 328 843
rect 341 839 346 843
rect 406 831 411 843
rect 424 839 429 843
rect 324 826 346 831
rect 406 826 429 831
rect 77 814 82 821
rect 93 814 98 821
rect 109 804 114 821
rect 125 804 130 821
rect 212 820 217 825
rect 272 820 277 825
rect 304 814 328 819
rect 304 806 309 814
rect 323 809 328 814
rect 341 809 346 826
rect 406 809 411 813
rect 424 809 429 826
rect 484 809 489 812
rect 323 786 328 804
rect 341 798 346 804
rect 406 786 411 804
rect 323 781 411 786
rect 424 769 429 804
rect 484 795 489 804
rect 485 791 489 795
rect 484 787 489 791
rect 484 777 489 782
rect 341 694 379 695
rect 384 694 429 695
rect 341 690 429 694
rect 212 677 217 680
rect 272 677 277 680
rect 323 673 328 677
rect 341 673 346 690
rect 406 673 411 677
rect 424 673 429 690
rect 212 663 217 672
rect 213 659 217 663
rect 212 655 217 659
rect 272 663 277 672
rect 272 659 276 663
rect 272 655 277 659
rect 323 656 328 668
rect 341 664 346 668
rect 406 656 411 668
rect 424 664 429 668
rect 324 651 346 656
rect 406 651 429 656
rect 212 645 217 650
rect 272 645 277 650
rect 304 639 328 644
rect 304 631 309 639
rect 323 634 328 639
rect 341 634 346 651
rect 406 634 411 638
rect 424 634 429 651
rect 484 634 489 637
rect 323 611 328 629
rect 341 623 346 629
rect 406 611 411 629
rect 323 606 411 611
rect 424 594 429 629
rect 484 620 489 629
rect 485 616 489 620
rect 484 612 489 616
rect 484 602 489 607
<< polycontact >>
rect 882 1562 887 1566
rect 936 1536 941 1542
rect 959 1536 964 1542
rect 774 1480 779 1484
rect 831 1481 836 1485
rect 669 1435 674 1442
rect 685 1435 690 1442
rect 701 1435 706 1442
rect 717 1436 722 1443
rect 722 1310 727 1315
rect 738 1310 744 1316
rect 883 1310 889 1317
rect 899 1310 905 1317
rect 931 1310 937 1316
rect 1060 1312 1067 1318
rect 379 1276 384 1281
rect 639 1277 644 1281
rect 1075 1310 1085 1318
rect 828 1277 833 1281
rect 986 1277 991 1281
rect 208 1241 213 1245
rect 1144 1259 1149 1263
rect 276 1241 281 1245
rect 319 1233 324 1238
rect 915 1229 922 1235
rect 1043 1229 1051 1236
rect 1198 1233 1203 1239
rect 1221 1233 1226 1239
rect 304 1208 309 1213
rect 480 1198 485 1202
rect 424 1171 429 1176
rect 376 1054 381 1059
rect 205 1019 210 1023
rect 273 1019 278 1023
rect 316 1011 321 1016
rect 301 986 306 991
rect 697 1013 702 1017
rect 844 1013 849 1017
rect 751 987 756 993
rect 774 987 779 993
rect 898 987 903 993
rect 990 1011 995 1015
rect 1126 1011 1131 1015
rect 921 987 926 993
rect 1044 985 1049 991
rect 1067 985 1072 991
rect 1180 985 1185 991
rect 1203 985 1208 991
rect 477 976 482 980
rect 421 949 426 954
rect 688 906 693 910
rect 833 905 838 909
rect 77 879 83 886
rect 93 879 99 886
rect 742 880 747 886
rect 765 880 770 886
rect 887 879 892 885
rect 982 903 987 907
rect 1126 903 1131 907
rect 910 879 915 885
rect 1036 877 1041 883
rect 1059 877 1064 883
rect 1180 877 1185 883
rect 1203 877 1208 883
rect 379 869 384 874
rect 22 846 27 850
rect 208 834 213 838
rect 276 834 281 838
rect 319 826 324 831
rect 109 798 116 804
rect 125 798 132 804
rect 304 801 309 806
rect 480 791 485 795
rect 424 764 429 769
rect 379 694 384 699
rect 208 659 213 663
rect 276 659 281 663
rect 319 651 324 656
rect 304 626 309 631
rect 480 616 485 620
rect 424 589 429 594
<< metal1 >>
rect 904 1606 932 1607
rect 904 1603 990 1606
rect 904 1593 908 1603
rect 929 1602 990 1603
rect 929 1601 980 1602
rect 929 1595 934 1601
rect 966 1595 971 1601
rect 904 1592 909 1593
rect 861 1587 909 1592
rect 975 1595 980 1601
rect 885 1580 890 1587
rect 897 1580 902 1587
rect 947 1580 952 1590
rect 947 1576 957 1580
rect 870 1566 875 1575
rect 953 1572 957 1576
rect 916 1569 957 1572
rect 916 1566 919 1569
rect 953 1566 957 1569
rect 859 1562 875 1566
rect 887 1562 919 1566
rect 870 1558 875 1562
rect 927 1561 929 1564
rect 885 1549 890 1553
rect 927 1550 930 1561
rect 944 1558 947 1561
rect 971 1550 974 1564
rect 859 1544 895 1549
rect 859 1543 866 1544
rect 927 1545 974 1550
rect 859 1522 864 1543
rect 936 1535 941 1536
rect 959 1520 964 1536
rect 950 1517 964 1520
rect 809 1510 857 1511
rect 985 1510 990 1602
rect 1247 1510 1270 1511
rect 647 1507 1271 1510
rect 647 1506 1262 1507
rect 647 1505 800 1506
rect 661 1494 666 1505
rect 737 1494 742 1505
rect 759 1498 764 1505
rect 771 1498 776 1505
rect 816 1499 821 1506
rect 828 1499 833 1506
rect 725 1467 730 1489
rect 786 1484 791 1493
rect 843 1485 848 1494
rect 944 1485 948 1493
rect 795 1484 831 1485
rect 756 1480 774 1484
rect 786 1481 831 1484
rect 843 1481 948 1485
rect 786 1480 829 1481
rect 756 1467 759 1480
rect 786 1476 791 1480
rect 843 1477 848 1481
rect 771 1467 776 1471
rect 828 1468 833 1472
rect 819 1467 858 1468
rect 677 1463 759 1467
rect 762 1463 882 1467
rect 677 1458 682 1463
rect 709 1458 714 1463
rect 762 1462 801 1463
rect 889 1463 1181 1467
rect 661 1449 666 1453
rect 693 1450 698 1453
rect 725 1450 730 1453
rect 762 1450 767 1462
rect 693 1449 767 1450
rect 661 1446 767 1449
rect 669 1433 674 1435
rect 685 1431 690 1435
rect 685 1418 689 1431
rect 701 1430 706 1435
rect 722 1436 866 1437
rect 717 1432 866 1436
rect 1178 1436 1181 1463
rect 1266 1454 1271 1507
rect 685 1415 795 1418
rect 292 1406 934 1408
rect 292 1405 935 1406
rect 292 1341 295 1405
rect 655 1382 660 1397
rect 796 1382 800 1397
rect 931 1384 935 1405
rect 141 1338 295 1341
rect 178 1337 295 1338
rect 578 1370 585 1373
rect 928 1370 952 1371
rect 578 1367 1066 1370
rect 94 1315 186 1317
rect 93 1310 186 1315
rect 76 887 82 1296
rect 77 886 82 887
rect 93 1077 99 1310
rect 460 1296 461 1302
rect 475 1296 554 1302
rect 379 1283 530 1288
rect 178 1279 372 1283
rect 178 1245 183 1279
rect 193 1267 356 1271
rect 193 1266 308 1267
rect 193 1259 198 1266
rect 205 1259 210 1266
rect 279 1259 284 1266
rect 220 1245 225 1254
rect 291 1259 296 1266
rect 303 1255 308 1266
rect 178 1242 208 1245
rect 204 1241 208 1242
rect 220 1241 229 1245
rect 264 1245 269 1254
rect 315 1255 320 1267
rect 238 1241 269 1245
rect 281 1241 287 1245
rect 220 1237 225 1241
rect 205 1228 210 1232
rect 196 1223 227 1228
rect 238 1177 242 1241
rect 264 1237 269 1241
rect 294 1241 302 1245
rect 298 1238 302 1241
rect 349 1244 354 1250
rect 367 1244 372 1279
rect 379 1281 384 1283
rect 398 1261 451 1267
rect 398 1255 403 1261
rect 432 1244 437 1250
rect 349 1239 437 1244
rect 298 1233 319 1238
rect 279 1228 284 1232
rect 255 1223 293 1228
rect 283 1186 288 1223
rect 349 1216 354 1239
rect 304 1205 309 1208
rect 383 1215 389 1228
rect 315 1186 320 1211
rect 398 1216 403 1226
rect 432 1216 437 1239
rect 446 1186 451 1261
rect 463 1223 506 1228
rect 465 1216 470 1223
rect 477 1216 482 1223
rect 492 1203 497 1211
rect 511 1203 516 1283
rect 548 1213 554 1296
rect 578 1248 585 1367
rect 717 1357 736 1362
rect 607 1231 611 1356
rect 655 1319 660 1356
rect 717 1321 725 1357
rect 796 1321 800 1359
rect 853 1327 889 1334
rect 717 1320 743 1321
rect 717 1318 744 1320
rect 736 1316 744 1318
rect 690 1310 722 1315
rect 736 1314 738 1316
rect 882 1318 888 1327
rect 883 1317 888 1318
rect 899 1317 904 1322
rect 931 1316 935 1358
rect 1061 1318 1066 1367
rect 1077 1336 1081 1386
rect 1178 1328 1182 1436
rect 1265 1434 1271 1454
rect 1077 1318 1081 1325
rect 617 1303 1130 1307
rect 1265 1305 1270 1434
rect 1248 1304 1306 1305
rect 618 1302 666 1303
rect 642 1295 647 1302
rect 654 1295 659 1302
rect 698 1291 703 1303
rect 730 1291 735 1303
rect 762 1291 767 1303
rect 807 1302 855 1303
rect 627 1281 632 1290
rect 831 1295 836 1302
rect 682 1283 687 1286
rect 714 1283 719 1286
rect 682 1282 719 1283
rect 746 1282 751 1286
rect 622 1277 632 1281
rect 644 1278 668 1281
rect 644 1277 659 1278
rect 627 1273 632 1277
rect 642 1264 647 1268
rect 664 1269 668 1278
rect 682 1278 751 1282
rect 796 1281 800 1291
rect 843 1295 848 1302
rect 863 1291 868 1303
rect 816 1281 821 1290
rect 875 1291 880 1303
rect 907 1291 912 1303
rect 939 1291 944 1303
rect 965 1302 1130 1303
rect 989 1295 994 1302
rect 1001 1295 1006 1302
rect 1027 1290 1032 1302
rect 1053 1290 1058 1302
rect 1085 1290 1090 1302
rect 891 1283 896 1286
rect 876 1282 896 1283
rect 923 1282 928 1286
rect 682 1269 687 1278
rect 796 1277 821 1281
rect 833 1277 852 1281
rect 664 1264 687 1269
rect 816 1273 821 1277
rect 831 1264 836 1268
rect 848 1269 852 1277
rect 876 1278 928 1282
rect 876 1269 881 1278
rect 974 1281 979 1290
rect 1036 1285 1037 1290
rect 1124 1289 1130 1302
rect 1163 1303 1194 1304
rect 1241 1303 1306 1304
rect 1163 1300 1306 1303
rect 1167 1289 1171 1300
rect 1036 1282 1042 1285
rect 1069 1282 1074 1285
rect 1123 1284 1171 1289
rect 1191 1298 1242 1300
rect 1248 1299 1306 1300
rect 1191 1292 1196 1298
rect 1228 1292 1233 1298
rect 1237 1292 1242 1298
rect 967 1277 979 1281
rect 991 1277 1017 1281
rect 1036 1277 1074 1282
rect 1147 1277 1152 1284
rect 848 1264 881 1269
rect 974 1273 979 1277
rect 989 1264 994 1268
rect 1013 1264 1017 1277
rect 1034 1264 1039 1277
rect 1159 1277 1164 1284
rect 1209 1277 1214 1287
rect 1209 1273 1219 1277
rect 617 1259 656 1264
rect 651 1243 656 1259
rect 682 1257 687 1264
rect 806 1259 845 1264
rect 762 1245 767 1252
rect 840 1245 845 1259
rect 876 1257 881 1264
rect 963 1259 1009 1264
rect 1013 1259 1039 1264
rect 762 1243 845 1245
rect 939 1250 944 1252
rect 964 1250 970 1259
rect 939 1247 970 1250
rect 1005 1258 1009 1259
rect 939 1246 949 1247
rect 939 1243 944 1246
rect 651 1240 944 1243
rect 1005 1244 1010 1258
rect 1034 1256 1039 1259
rect 1132 1263 1137 1272
rect 1215 1269 1219 1273
rect 1178 1266 1219 1269
rect 1178 1263 1181 1266
rect 1215 1263 1219 1266
rect 1126 1259 1137 1263
rect 1149 1259 1181 1263
rect 1085 1244 1090 1251
rect 1132 1255 1137 1259
rect 1189 1258 1191 1261
rect 1147 1246 1152 1250
rect 1189 1247 1192 1258
rect 1206 1255 1209 1258
rect 1233 1247 1236 1261
rect 1121 1244 1157 1246
rect 1005 1241 1157 1244
rect 1005 1240 1130 1241
rect 1189 1242 1236 1247
rect 651 1239 767 1240
rect 840 1239 944 1240
rect 607 1229 690 1231
rect 607 1227 695 1229
rect 706 1222 711 1229
rect 754 1226 759 1229
rect 706 1218 737 1222
rect 548 1211 683 1213
rect 548 1208 684 1211
rect 477 1198 480 1202
rect 492 1198 516 1203
rect 492 1194 497 1198
rect 678 1194 684 1208
rect 728 1207 736 1218
rect 730 1199 736 1207
rect 753 1213 762 1226
rect 915 1225 920 1229
rect 1045 1226 1049 1229
rect 753 1206 755 1213
rect 728 1198 736 1199
rect 283 1185 451 1186
rect 477 1185 482 1189
rect 283 1181 530 1185
rect 446 1180 530 1181
rect 238 1172 407 1177
rect 402 1167 407 1172
rect 424 1167 429 1171
rect 402 1162 429 1167
rect 93 1074 224 1077
rect 93 1073 99 1074
rect 93 886 98 1073
rect 507 1066 514 1132
rect 376 1061 514 1066
rect 175 1057 369 1061
rect 175 1023 180 1057
rect 190 1045 353 1049
rect 190 1044 305 1045
rect 190 1037 195 1044
rect 202 1037 207 1044
rect 276 1037 281 1044
rect 217 1023 222 1032
rect 288 1037 293 1044
rect 300 1033 305 1044
rect 175 1020 205 1023
rect 201 1019 205 1020
rect 217 1019 226 1023
rect 261 1023 266 1032
rect 312 1033 317 1045
rect 235 1019 266 1023
rect 278 1021 299 1023
rect 278 1019 286 1021
rect 217 1015 222 1019
rect 202 1006 207 1010
rect 193 1001 224 1006
rect 235 955 239 1019
rect 261 1015 266 1019
rect 292 1019 299 1021
rect 295 1016 299 1019
rect 346 1022 351 1028
rect 364 1022 369 1057
rect 376 1059 381 1061
rect 395 1039 448 1045
rect 395 1033 400 1039
rect 429 1022 434 1028
rect 346 1017 434 1022
rect 295 1011 316 1016
rect 276 1006 281 1010
rect 252 1001 290 1006
rect 280 964 285 1001
rect 346 994 351 1017
rect 395 1011 398 1014
rect 388 1006 403 1011
rect 301 983 306 986
rect 380 995 385 1006
rect 395 994 400 1006
rect 429 994 434 1017
rect 312 964 317 989
rect 443 964 448 1039
rect 460 1001 503 1006
rect 462 994 467 1001
rect 474 994 479 1001
rect 489 981 494 989
rect 508 981 513 1061
rect 474 976 477 980
rect 489 976 513 981
rect 523 998 529 1180
rect 548 1143 557 1181
rect 677 1188 684 1194
rect 570 1129 577 1180
rect 620 1156 621 1163
rect 620 1099 627 1156
rect 552 1091 628 1099
rect 677 1091 683 1188
rect 739 1150 748 1175
rect 914 1171 920 1225
rect 1044 1163 1049 1226
rect 1121 1218 1130 1240
rect 1198 1232 1203 1233
rect 1221 1232 1226 1233
rect 1122 1209 1130 1218
rect 1122 1206 1306 1209
rect 739 1144 1109 1150
rect 789 1112 815 1118
rect 1102 1110 1109 1144
rect 727 1095 958 1099
rect 676 1086 683 1091
rect 585 1065 651 1072
rect 677 1043 683 1086
rect 716 1057 747 1058
rect 794 1057 894 1058
rect 716 1056 942 1057
rect 716 1055 1040 1056
rect 1145 1055 1176 1056
rect 716 1054 1306 1055
rect 720 1043 724 1054
rect 676 1038 724 1043
rect 744 1052 795 1054
rect 744 1046 749 1052
rect 781 1046 786 1052
rect 790 1046 795 1052
rect 867 1043 871 1054
rect 700 1031 705 1038
rect 712 1031 717 1038
rect 762 1031 767 1041
rect 823 1038 871 1043
rect 891 1052 1306 1054
rect 891 1046 896 1052
rect 928 1046 933 1052
rect 937 1046 942 1052
rect 1013 1041 1017 1052
rect 847 1031 852 1038
rect 762 1027 772 1031
rect 685 1017 690 1026
rect 768 1023 772 1027
rect 731 1020 772 1023
rect 731 1017 734 1020
rect 768 1017 772 1020
rect 859 1031 864 1038
rect 909 1031 914 1041
rect 969 1036 1017 1041
rect 1037 1051 1153 1052
rect 1037 1050 1088 1051
rect 1037 1044 1042 1050
rect 1074 1044 1079 1050
rect 1083 1044 1088 1050
rect 1149 1041 1153 1051
rect 909 1027 919 1031
rect 993 1029 998 1036
rect 667 1013 690 1017
rect 702 1013 734 1017
rect 685 1009 690 1013
rect 742 1012 744 1015
rect 700 1000 705 1004
rect 742 1001 745 1012
rect 759 1009 762 1012
rect 786 1001 789 1015
rect 832 1017 837 1026
rect 915 1023 919 1027
rect 878 1020 919 1023
rect 878 1017 881 1020
rect 915 1017 919 1020
rect 1005 1029 1010 1036
rect 1055 1029 1060 1039
rect 1105 1036 1153 1041
rect 1173 1050 1306 1052
rect 1173 1044 1178 1050
rect 1210 1044 1215 1050
rect 1218 1049 1306 1050
rect 1219 1044 1224 1049
rect 1129 1029 1134 1036
rect 1055 1025 1065 1029
rect 821 1014 837 1017
rect 819 1013 837 1014
rect 849 1013 881 1017
rect 832 1009 837 1013
rect 889 1012 891 1015
rect 674 998 710 1000
rect 523 995 710 998
rect 523 993 683 995
rect 742 996 789 1001
rect 847 1000 852 1004
rect 889 1001 892 1012
rect 906 1009 909 1012
rect 933 1001 936 1015
rect 978 1015 983 1024
rect 1061 1021 1065 1025
rect 1024 1018 1065 1021
rect 1024 1015 1027 1018
rect 1061 1015 1065 1018
rect 1141 1029 1146 1036
rect 1191 1029 1196 1039
rect 1191 1025 1201 1029
rect 1114 1015 1119 1024
rect 1197 1021 1201 1025
rect 1160 1018 1201 1021
rect 1160 1015 1163 1018
rect 1197 1015 1201 1018
rect 966 1011 983 1015
rect 995 1011 1027 1015
rect 978 1007 983 1011
rect 1035 1010 1037 1013
rect 1104 1014 1119 1015
rect 819 995 857 1000
rect 489 972 494 976
rect 280 963 448 964
rect 474 963 479 967
rect 523 963 529 993
rect 280 959 529 963
rect 443 958 529 959
rect 235 950 404 955
rect 399 945 404 950
rect 421 945 426 949
rect 160 934 198 938
rect 399 940 426 945
rect 160 933 202 934
rect 483 881 488 893
rect 144 876 149 881
rect 379 876 516 881
rect 1 872 149 876
rect 153 872 372 876
rect 1 871 49 872
rect 25 864 30 871
rect 37 864 42 871
rect 57 860 62 872
rect 10 850 15 859
rect 69 860 74 872
rect 101 860 106 872
rect 133 860 138 872
rect 85 852 90 855
rect 70 851 90 852
rect 117 851 122 855
rect 3 846 15 850
rect 27 846 46 850
rect 10 842 15 846
rect 25 833 30 837
rect 42 838 46 846
rect 70 847 122 851
rect 70 838 75 847
rect 42 833 45 838
rect 50 833 75 838
rect 153 838 158 872
rect 168 860 356 864
rect 168 859 308 860
rect 168 852 173 859
rect 205 852 210 859
rect 279 852 284 859
rect 220 838 225 847
rect 291 852 296 859
rect 303 848 308 859
rect 264 838 269 847
rect 315 848 320 860
rect 153 835 208 838
rect 204 834 208 835
rect 220 834 228 838
rect 0 828 39 833
rect 34 812 39 828
rect 70 826 75 833
rect 220 830 225 834
rect 238 834 269 838
rect 281 836 302 838
rect 281 834 288 836
rect 205 821 210 825
rect 133 819 138 821
rect 171 819 227 821
rect 133 816 227 819
rect 133 815 175 816
rect 133 812 138 815
rect 34 808 138 812
rect 153 801 186 804
rect 109 782 114 798
rect 125 793 130 798
rect 125 789 226 793
rect 109 778 143 782
rect 238 770 242 834
rect 264 830 269 834
rect 293 834 302 836
rect 298 831 302 834
rect 349 837 354 843
rect 367 837 372 872
rect 379 874 384 876
rect 398 854 451 860
rect 398 848 403 854
rect 432 837 437 843
rect 349 832 437 837
rect 298 826 319 831
rect 279 821 284 825
rect 255 816 293 821
rect 283 779 288 816
rect 349 809 354 832
rect 398 826 401 829
rect 304 798 309 801
rect 391 821 406 826
rect 383 808 388 821
rect 315 779 320 804
rect 398 809 403 821
rect 432 809 437 832
rect 446 779 451 854
rect 463 816 506 821
rect 465 809 470 816
rect 477 809 482 816
rect 492 796 497 804
rect 511 796 516 876
rect 477 791 480 795
rect 492 791 516 796
rect 492 787 497 791
rect 283 778 451 779
rect 477 778 482 782
rect 523 778 529 958
rect 541 965 542 974
rect 647 972 655 973
rect 674 972 683 993
rect 751 986 756 987
rect 774 986 779 987
rect 819 972 828 995
rect 889 996 936 1001
rect 993 998 998 1002
rect 1035 999 1038 1010
rect 1052 1007 1055 1010
rect 1079 999 1082 1013
rect 1109 1011 1119 1014
rect 1131 1011 1163 1015
rect 1114 1007 1119 1011
rect 1171 1010 1173 1013
rect 968 997 1003 998
rect 955 993 1003 997
rect 898 986 903 987
rect 955 992 974 993
rect 1035 994 1082 999
rect 1129 998 1134 1002
rect 1171 999 1174 1010
rect 1188 1007 1191 1010
rect 1215 999 1218 1013
rect 1104 993 1139 998
rect 921 986 926 987
rect 957 972 964 992
rect 1044 984 1049 985
rect 1067 984 1072 985
rect 1104 972 1108 993
rect 1171 994 1218 999
rect 1180 984 1185 985
rect 1203 984 1208 985
rect 541 922 548 965
rect 575 888 581 971
rect 647 966 1108 972
rect 545 882 581 888
rect 618 857 620 866
rect 618 789 627 857
rect 283 774 531 778
rect 446 773 531 774
rect 238 765 407 770
rect 402 760 407 765
rect 424 760 429 764
rect 402 755 429 760
rect 502 736 506 758
rect 379 701 510 706
rect 178 697 372 701
rect 178 663 183 697
rect 193 685 356 689
rect 193 684 308 685
rect 193 677 198 684
rect 205 677 210 684
rect 279 677 284 684
rect 220 663 225 672
rect 291 677 296 684
rect 303 673 308 684
rect 264 663 269 672
rect 315 673 320 685
rect 178 660 208 663
rect 204 659 208 660
rect 220 659 228 663
rect 220 655 225 659
rect 238 659 269 663
rect 281 661 302 663
rect 281 659 288 661
rect 205 646 210 650
rect 196 641 227 646
rect 238 595 242 659
rect 264 655 269 659
rect 294 659 302 661
rect 298 656 302 659
rect 349 662 354 668
rect 367 662 372 697
rect 379 699 384 701
rect 398 679 451 685
rect 398 673 403 679
rect 432 662 437 668
rect 349 657 437 662
rect 298 651 319 656
rect 279 646 284 650
rect 255 641 293 646
rect 283 604 288 641
rect 349 634 354 657
rect 398 651 401 654
rect 388 646 406 651
rect 304 623 309 626
rect 379 634 386 646
rect 398 634 403 646
rect 379 629 383 634
rect 432 634 437 657
rect 315 604 320 629
rect 446 604 451 679
rect 463 641 506 646
rect 465 634 470 641
rect 477 634 482 641
rect 492 621 497 629
rect 511 621 516 701
rect 477 616 480 620
rect 492 616 516 621
rect 492 612 497 616
rect 283 603 451 604
rect 477 603 482 607
rect 523 603 529 773
rect 617 705 627 789
rect 617 640 626 705
rect 283 599 529 603
rect 446 598 529 599
rect 238 590 407 595
rect 402 585 407 590
rect 424 585 429 589
rect 402 580 429 585
rect 476 562 483 571
rect 635 562 641 906
rect 647 860 655 966
rect 707 950 738 951
rect 707 949 883 950
rect 1237 949 1245 1049
rect 707 948 1007 949
rect 707 947 1032 948
rect 1145 947 1176 948
rect 1215 947 1245 949
rect 711 936 715 947
rect 667 931 715 936
rect 735 946 1245 947
rect 735 945 871 946
rect 735 939 740 945
rect 772 939 777 945
rect 781 939 786 945
rect 856 935 860 945
rect 691 924 696 931
rect 703 924 708 931
rect 753 924 758 934
rect 812 930 860 935
rect 880 944 1245 946
rect 880 938 885 944
rect 917 938 922 944
rect 926 938 931 944
rect 1005 933 1009 944
rect 753 920 763 924
rect 836 923 841 930
rect 676 910 681 919
rect 759 916 763 920
rect 722 913 763 916
rect 722 910 725 913
rect 759 910 763 913
rect 848 923 853 930
rect 898 923 903 933
rect 961 928 1009 933
rect 1029 942 1154 944
rect 1173 942 1245 944
rect 1029 936 1034 942
rect 1066 936 1071 942
rect 1075 936 1080 942
rect 1149 933 1153 942
rect 898 919 908 923
rect 985 921 990 928
rect 668 906 681 910
rect 693 906 725 910
rect 676 902 681 906
rect 733 905 735 908
rect 665 893 672 894
rect 691 893 696 897
rect 733 894 736 905
rect 750 902 753 905
rect 777 894 780 908
rect 821 909 826 918
rect 904 915 908 919
rect 867 912 908 915
rect 867 909 870 912
rect 904 909 908 912
rect 997 921 1002 928
rect 1047 921 1052 931
rect 1105 928 1153 933
rect 1173 936 1178 942
rect 1210 936 1215 942
rect 1219 936 1224 942
rect 1129 921 1134 928
rect 1047 917 1057 921
rect 809 906 826 909
rect 818 905 826 906
rect 838 905 870 909
rect 821 901 826 905
rect 878 904 880 907
rect 970 907 975 916
rect 1053 913 1057 917
rect 1016 910 1057 913
rect 1016 907 1019 910
rect 1053 907 1057 910
rect 1141 921 1146 928
rect 1191 921 1196 931
rect 1191 917 1201 921
rect 665 888 701 893
rect 665 861 672 888
rect 733 889 780 894
rect 836 892 841 896
rect 878 893 881 904
rect 895 901 898 904
rect 922 893 925 907
rect 952 902 975 907
rect 987 903 1019 907
rect 970 899 975 902
rect 1027 902 1029 905
rect 811 887 846 892
rect 742 879 747 880
rect 765 878 770 880
rect 811 861 818 887
rect 878 888 925 893
rect 985 890 990 894
rect 1027 891 1030 902
rect 1044 899 1047 902
rect 1071 891 1074 905
rect 1114 907 1119 916
rect 1197 913 1201 917
rect 1160 910 1201 913
rect 1160 907 1163 910
rect 1197 907 1201 910
rect 1095 903 1119 907
rect 1131 903 1163 907
rect 1114 899 1119 903
rect 1171 902 1173 905
rect 954 885 995 890
rect 887 878 892 879
rect 910 878 915 879
rect 955 861 962 885
rect 1027 886 1074 891
rect 1129 890 1134 894
rect 1171 891 1174 902
rect 1188 899 1191 902
rect 1215 891 1218 905
rect 1104 885 1139 890
rect 1036 876 1041 877
rect 1059 876 1064 877
rect 1103 861 1112 885
rect 1171 886 1218 891
rect 1180 876 1185 877
rect 1203 876 1208 877
rect 1249 868 1306 872
rect 665 860 1112 861
rect 647 855 1112 860
rect 665 854 672 855
rect 955 853 962 855
rect 1103 836 1111 855
rect 1103 832 1306 836
rect 476 556 641 562
rect 673 539 682 625
rect 299 533 682 539
<< m2contact >>
rect 944 1553 949 1558
rect 895 1543 902 1550
rect 936 1528 941 1535
rect 859 1517 869 1522
rect 944 1517 950 1522
rect 943 1493 949 1499
rect 882 1462 889 1469
rect 669 1426 674 1433
rect 866 1430 872 1439
rect 700 1424 707 1430
rect 795 1413 800 1419
rect 132 1335 141 1346
rect 655 1397 661 1402
rect 795 1397 802 1402
rect 1071 1386 1086 1395
rect 655 1377 662 1382
rect 795 1377 802 1382
rect 931 1379 936 1384
rect 186 1310 199 1320
rect 75 1296 86 1306
rect 461 1294 475 1304
rect 186 1266 193 1272
rect 229 1241 234 1246
rect 356 1266 361 1271
rect 227 1223 232 1228
rect 287 1240 294 1245
rect 250 1223 255 1228
rect 304 1200 309 1205
rect 383 1228 390 1235
rect 398 1226 403 1233
rect 458 1223 463 1228
rect 530 1282 538 1290
rect 604 1356 615 1363
rect 655 1356 663 1362
rect 736 1357 750 1362
rect 795 1359 802 1364
rect 578 1234 587 1248
rect 931 1358 937 1363
rect 840 1322 853 1338
rect 655 1312 664 1319
rect 681 1310 690 1318
rect 796 1315 801 1321
rect 899 1322 909 1331
rect 1077 1325 1088 1336
rect 1176 1319 1187 1328
rect 796 1291 801 1298
rect 615 1276 622 1281
rect 961 1275 967 1283
rect 1116 1258 1126 1264
rect 1206 1250 1211 1255
rect 1157 1240 1164 1247
rect 690 1229 695 1235
rect 706 1229 711 1235
rect 754 1229 759 1236
rect 472 1198 477 1203
rect 720 1199 730 1207
rect 755 1205 765 1213
rect 545 1181 561 1193
rect 503 1132 517 1141
rect 224 1072 229 1077
rect 183 1043 190 1049
rect 226 1019 231 1024
rect 353 1044 358 1049
rect 224 1001 229 1006
rect 286 1015 292 1021
rect 247 1001 252 1006
rect 379 1006 388 1011
rect 301 978 306 983
rect 455 1001 460 1006
rect 469 976 474 981
rect 568 1180 585 1191
rect 548 1131 560 1143
rect 621 1156 633 1167
rect 570 1114 581 1129
rect 541 1091 552 1102
rect 739 1175 751 1191
rect 914 1162 925 1171
rect 1198 1225 1203 1232
rect 1221 1225 1226 1232
rect 1012 1156 1024 1163
rect 1039 1156 1051 1163
rect 779 1112 789 1119
rect 815 1110 828 1120
rect 716 1095 727 1106
rect 958 1093 970 1107
rect 1102 1101 1117 1110
rect 573 1064 585 1074
rect 651 1065 662 1074
rect 660 1013 667 1019
rect 759 1004 764 1009
rect 815 1014 821 1019
rect 710 994 717 1001
rect 906 1004 911 1009
rect 959 1011 966 1017
rect 153 933 160 940
rect 198 934 205 941
rect 480 893 489 903
rect 144 881 152 887
rect 45 833 50 838
rect 161 859 168 865
rect 356 859 361 864
rect 228 832 233 838
rect 227 816 232 821
rect 147 800 153 806
rect 186 800 192 805
rect 226 788 231 794
rect 143 776 151 782
rect 288 831 293 836
rect 250 816 255 821
rect 304 793 309 798
rect 383 821 391 826
rect 458 816 463 821
rect 472 791 477 796
rect 542 965 554 976
rect 572 971 583 981
rect 751 979 756 986
rect 774 979 779 986
rect 857 994 864 1001
rect 1052 1002 1057 1007
rect 1103 1009 1109 1014
rect 898 979 903 986
rect 1003 992 1010 999
rect 1188 1002 1193 1007
rect 921 979 926 986
rect 1044 977 1049 984
rect 1067 977 1072 984
rect 1139 992 1146 999
rect 1180 977 1185 984
rect 1203 977 1208 984
rect 541 909 551 922
rect 535 882 545 890
rect 635 906 641 911
rect 620 857 630 867
rect 501 758 510 765
rect 502 729 509 736
rect 510 701 516 709
rect 186 684 193 690
rect 356 684 361 689
rect 228 658 233 663
rect 227 641 232 646
rect 288 656 294 661
rect 250 641 255 646
rect 378 646 388 651
rect 304 618 309 623
rect 458 641 463 646
rect 472 616 477 621
rect 617 628 626 640
rect 476 571 485 581
rect 662 904 668 910
rect 750 897 755 902
rect 804 906 809 911
rect 701 887 708 894
rect 895 896 900 901
rect 945 902 952 907
rect 742 872 747 879
rect 765 871 770 878
rect 846 886 853 893
rect 1044 894 1049 899
rect 1090 903 1095 908
rect 887 871 892 878
rect 910 871 915 878
rect 995 884 1002 891
rect 1188 894 1193 899
rect 1036 869 1041 876
rect 1059 869 1064 876
rect 1139 884 1146 891
rect 1180 869 1185 876
rect 1203 868 1208 876
rect 1244 868 1249 874
rect 671 625 685 640
rect 288 533 299 544
<< metal2 >>
rect 918 1553 944 1556
rect 918 1549 923 1553
rect 902 1544 923 1549
rect 632 1528 936 1531
rect 632 1526 941 1528
rect 633 1447 636 1526
rect 869 1517 888 1522
rect 883 1469 888 1517
rect 944 1499 947 1517
rect 46 1444 636 1447
rect 46 1294 50 1444
rect 655 1426 669 1428
rect 872 1432 906 1437
rect 655 1424 674 1426
rect 707 1425 824 1428
rect 754 1424 824 1425
rect 655 1402 659 1424
rect 796 1402 800 1413
rect 342 1389 1071 1393
rect 125 1337 132 1342
rect 343 1321 348 1389
rect 554 1358 604 1362
rect 655 1362 660 1377
rect 742 1362 746 1389
rect 796 1364 800 1377
rect 931 1363 935 1379
rect 571 1348 1257 1352
rect 199 1310 283 1318
rect 178 1302 234 1303
rect 86 1300 234 1302
rect 343 1300 349 1321
rect 86 1297 349 1300
rect 86 1296 184 1297
rect 45 1213 50 1294
rect 45 838 49 1213
rect 154 940 158 1273
rect 186 1049 189 1266
rect 229 1246 234 1297
rect 364 1294 461 1300
rect 364 1291 471 1294
rect 364 1271 369 1291
rect 361 1266 383 1271
rect 232 1223 250 1228
rect 288 1123 293 1240
rect 377 1228 383 1266
rect 390 1228 398 1233
rect 458 1228 463 1291
rect 571 1287 580 1348
rect 731 1331 840 1332
rect 645 1326 840 1331
rect 645 1325 759 1326
rect 538 1282 580 1287
rect 615 1312 655 1317
rect 681 1318 688 1325
rect 853 1326 856 1332
rect 1008 1327 1077 1330
rect 909 1325 1077 1327
rect 909 1322 1081 1325
rect 615 1281 621 1312
rect 796 1298 800 1315
rect 961 1283 966 1311
rect 1116 1264 1120 1325
rect 1177 1253 1182 1319
rect 1251 1307 1257 1348
rect 1177 1250 1206 1253
rect 556 1239 578 1245
rect 304 1158 309 1200
rect 462 1198 472 1202
rect 462 1158 468 1198
rect 556 1193 562 1239
rect 1177 1246 1185 1250
rect 1164 1241 1185 1246
rect 1250 1230 1257 1307
rect 1226 1227 1257 1230
rect 1226 1226 1254 1227
rect 1198 1221 1203 1225
rect 714 1199 720 1205
rect 561 1181 562 1193
rect 585 1180 739 1188
rect 304 1157 610 1158
rect 304 1153 612 1157
rect 633 1162 720 1163
rect 633 1156 721 1162
rect 457 1152 612 1153
rect 596 1150 612 1152
rect 517 1132 548 1139
rect 288 1118 570 1123
rect 186 892 189 1043
rect 226 1024 229 1072
rect 361 1069 468 1078
rect 361 1049 366 1069
rect 358 1044 380 1049
rect 229 1001 247 1006
rect 205 935 232 939
rect 161 888 189 892
rect 161 887 164 888
rect 152 881 164 887
rect 228 885 232 935
rect 287 916 291 1015
rect 374 1011 380 1044
rect 374 1006 379 1011
rect 455 1006 460 1069
rect 301 936 306 978
rect 459 976 469 980
rect 542 976 548 1091
rect 575 981 580 1064
rect 459 936 465 976
rect 301 933 465 936
rect 301 931 565 933
rect 454 930 565 931
rect 287 912 541 916
rect 398 897 480 901
rect 161 865 164 881
rect 200 882 232 885
rect 200 870 205 882
rect 186 867 205 870
rect 146 800 147 805
rect 146 782 149 800
rect 161 782 164 859
rect 186 805 190 867
rect 228 838 232 882
rect 364 884 471 893
rect 364 864 369 884
rect 361 859 383 864
rect 232 816 250 821
rect 161 778 189 782
rect 186 690 189 778
rect 228 663 231 788
rect 289 733 293 831
rect 377 821 383 859
rect 458 821 463 884
rect 304 751 309 793
rect 462 791 472 795
rect 462 751 468 791
rect 537 763 542 882
rect 560 861 565 930
rect 510 760 542 763
rect 510 759 541 760
rect 304 749 468 751
rect 558 750 565 861
rect 600 823 610 1150
rect 634 1124 640 1125
rect 634 1119 706 1124
rect 634 1021 640 1119
rect 699 1090 705 1119
rect 716 1106 721 1156
rect 758 1090 763 1205
rect 802 1185 1306 1195
rect 781 1096 787 1112
rect 699 1086 763 1090
rect 780 1072 787 1096
rect 662 1065 787 1072
rect 620 1020 656 1021
rect 620 1019 664 1020
rect 620 1015 660 1019
rect 620 867 628 1015
rect 633 1014 660 1015
rect 733 1004 759 1007
rect 733 1000 738 1004
rect 717 995 738 1000
rect 803 984 810 1185
rect 943 1167 1306 1174
rect 815 1088 819 1110
rect 918 1088 923 1162
rect 815 1084 924 1088
rect 815 1019 819 1084
rect 880 1004 906 1007
rect 880 1000 885 1004
rect 864 995 885 1000
rect 779 981 810 984
rect 779 980 807 981
rect 751 961 756 979
rect 898 961 903 979
rect 943 983 950 1167
rect 1007 1156 1012 1162
rect 1024 1156 1039 1163
rect 959 1087 963 1093
rect 1007 1087 1014 1156
rect 1092 1137 1306 1145
rect 959 1081 1015 1087
rect 959 1017 963 1081
rect 1026 1002 1052 1005
rect 1026 998 1031 1002
rect 1010 993 1031 998
rect 926 979 950 983
rect 921 978 948 979
rect 1092 980 1097 1137
rect 1253 1123 1260 1124
rect 1253 1117 1306 1123
rect 1103 1096 1109 1101
rect 1103 1090 1199 1096
rect 1103 1014 1109 1090
rect 1162 1002 1188 1005
rect 1162 998 1167 1002
rect 1146 993 1167 998
rect 1072 977 1098 980
rect 1044 961 1049 977
rect 1180 961 1185 977
rect 1253 979 1260 1117
rect 1208 977 1260 979
rect 1203 974 1260 977
rect 751 958 1270 961
rect 641 906 662 910
rect 724 897 750 900
rect 804 901 807 906
rect 724 893 729 897
rect 869 896 895 899
rect 708 888 729 893
rect 869 892 874 896
rect 853 887 874 892
rect 945 894 948 902
rect 1018 894 1044 897
rect 1018 890 1023 894
rect 1002 885 1023 890
rect 1090 883 1094 903
rect 1162 894 1188 897
rect 1162 890 1167 894
rect 1146 885 1167 890
rect 742 847 747 872
rect 770 872 792 876
rect 887 847 892 871
rect 915 871 931 873
rect 910 869 931 871
rect 1064 869 1074 873
rect 1036 847 1041 869
rect 1180 847 1185 869
rect 1208 868 1244 872
rect 1266 847 1270 958
rect 742 844 1270 847
rect 742 843 747 844
rect 600 820 1090 823
rect 600 819 610 820
rect 1266 814 1270 844
rect 896 799 900 804
rect 895 796 946 799
rect 953 796 954 799
rect 895 795 954 796
rect 772 781 805 784
rect 772 780 810 781
rect 558 749 616 750
rect 896 749 900 795
rect 1080 765 1162 771
rect 304 746 551 749
rect 289 729 502 733
rect 364 709 471 718
rect 510 709 516 715
rect 364 689 369 709
rect 361 684 383 689
rect 232 641 250 646
rect 288 561 292 656
rect 377 651 383 684
rect 377 646 378 651
rect 458 646 463 709
rect 304 576 309 618
rect 462 616 472 620
rect 462 577 468 616
rect 461 576 476 577
rect 304 571 476 576
rect 542 575 551 746
rect 558 746 903 749
rect 558 743 616 746
rect 940 745 1162 751
rect 800 717 1162 721
rect 626 628 671 637
rect 749 577 759 578
rect 631 576 759 577
rect 571 575 759 576
rect 542 572 759 575
rect 542 571 749 572
rect 288 544 293 561
<< m3contact >>
rect 906 1431 913 1437
rect 824 1421 837 1429
rect 113 1334 125 1346
rect 546 1357 554 1366
rect 283 1309 299 1321
rect 152 1273 160 1281
rect 631 1323 645 1334
rect 1114 1325 1127 1332
rect 959 1311 967 1316
rect 1197 1215 1205 1221
rect 706 1199 714 1207
rect 387 897 398 905
rect 1199 1090 1207 1096
rect 804 896 809 901
rect 945 889 950 894
rect 1090 878 1095 883
rect 792 872 797 878
rect 931 868 938 874
rect 1074 869 1080 876
rect 1090 819 1095 824
rect 946 796 953 802
rect 763 779 772 787
rect 805 781 812 787
rect 1072 765 1080 775
rect 510 715 517 723
rect 931 745 940 754
rect 795 717 800 725
rect 759 569 771 582
<< metal3 >>
rect 913 1431 1033 1436
rect 1029 1422 1033 1431
rect 829 1419 1000 1421
rect 1029 1419 1119 1422
rect 829 1417 1001 1419
rect 1029 1417 1121 1419
rect 154 1364 157 1365
rect 152 1359 546 1364
rect 116 926 120 1334
rect 154 1281 157 1359
rect 390 1330 394 1332
rect 535 1330 631 1331
rect 389 1326 631 1330
rect 390 1318 394 1326
rect 535 1324 631 1326
rect 299 1309 395 1318
rect 997 1316 1001 1417
rect 1116 1332 1121 1417
rect 967 1311 1002 1316
rect 607 1134 615 1136
rect 707 1134 712 1199
rect 606 1127 713 1134
rect 580 943 587 945
rect 607 943 615 1127
rect 1199 1096 1202 1215
rect 580 936 616 943
rect 116 922 248 926
rect 240 902 245 922
rect 240 898 387 902
rect 580 825 587 936
rect 797 872 798 877
rect 579 721 587 825
rect 517 715 587 721
rect 761 779 763 785
rect 761 582 766 779
rect 795 725 798 872
rect 806 787 809 896
rect 931 754 937 868
rect 946 802 949 889
rect 1073 869 1074 871
rect 1073 775 1079 869
rect 1090 824 1094 878
<< labels >>
rlabel metal1 1197 997 1197 997 1 compare_node_1
rlabel metal1 1058 997 1058 997 1 compare_node_2
rlabel metal1 912 998 912 998 1 compare_node_3
rlabel metal1 766 998 766 998 1 compare_node_4
rlabel metal1 757 892 757 892 1 compare_node_5
rlabel metal1 901 890 901 890 1 compare_node_6
rlabel metal1 1051 887 1051 887 1 compare_node_7
rlabel metal1 1194 887 1194 887 1 compare_node_8
rlabel metal1 1197 1028 1197 1028 1 compare_A3e_nand
rlabel metal1 1063 1027 1063 1027 1 compare_A2e_nand
rlabel metal1 917 1026 917 1026 1 compare_A1e_nand
rlabel metal1 769 1030 769 1030 1 compare_A0e_nand
rlabel metal1 761 923 761 923 1 compare_B0e_nand
rlabel metal1 906 920 906 920 1 compare_B1e_nand
rlabel metal1 1054 919 1054 919 1 compare_B2e_nand
rlabel metal1 1199 919 1199 919 1 compare_B3e_nand
rlabel metal1 1113 1013 1113 1013 1 compare_A3e
rlabel metal1 978 1014 978 1014 1 compare_A2e
rlabel metal1 834 1014 834 1014 1 compare_A1e
rlabel metal1 685 1016 685 1016 1 compare_A0e
rlabel metal1 677 908 677 908 1 compare_B0e
rlabel metal1 823 907 823 907 1 compare_B1e
rlabel metal1 972 904 972 904 1 compare_B2e
rlabel metal1 1117 905 1117 905 1 compare_B3e
rlabel pdiffusion 335 1253 335 1253 1 xnor_1
rlabel ndiffusion 335 1213 335 1213 1 xnor_2
rlabel metal1 396 1242 396 1242 1 xor_1
rlabel ndiffusion 417 1253 417 1253 1 xnor_3
rlabel pdiffusion 417 1213 417 1213 1 xnor_4
rlabel metal1 425 1167 425 1167 1 A3c
rlabel metal1 382 1284 382 1284 1 B3c
rlabel pdiffusion 330 1031 330 1031 1 xnor_5
rlabel ndiffusion 333 991 333 991 1 xnor_6
rlabel ndiffusion 416 1031 416 1031 1 xnor_7
rlabel pdiffusion 412 990 412 990 1 xnor_8
rlabel metal1 424 942 424 942 1 A2c
rlabel metal1 383 1064 383 1064 1 B2c
rlabel metal1 383 879 383 879 1 B1c
rlabel metal1 417 756 417 756 1 A1c
rlabel pdiffusion 335 845 335 845 1 xnor_9
rlabel ndiffusion 338 806 338 806 1 xnor_10
rlabel pdiffusion 416 806 416 806 1 xnor_11
rlabel ndiffusion 418 846 418 846 1 xnor_12
rlabel metal1 385 1018 385 1018 1 xor_2
rlabel metal1 390 834 390 834 1 xor_3
rlabel metal1 393 703 393 703 1 B0c
rlabel metal1 417 582 417 582 1 A0c
rlabel metal1 393 660 393 660 1 xor_4
rlabel pdiffusion 334 671 334 671 1 xnor_13
rlabel ndiffusion 336 630 336 630 1 xnor_14
rlabel ndiffusion 418 670 418 670 1 xnor_15
rlabel pdiffusion 418 631 418 631 1 xnor_16
rlabel ndiffusion 88 823 88 823 1 A_compare_B_node_3
rlabel ndiffusion 105 824 105 824 1 A_compare_B_node_2
rlabel ndiffusion 120 824 120 824 1 A_compare_B_node_1
rlabel metal1 5 848 5 848 3 A_equal_B
rlabel metal1 51 836 51 836 1 A_equal_B_c
rlabel metal1 94 906 94 906 1 A2e_xnor_B2e
rlabel metal1 223 1244 223 1244 1 A3e_xnor_B3e
rlabel metal1 222 836 222 836 1 A1e_xnor_B1e
rlabel metal1 223 660 223 660 1 A0e_xnor_B0e
rlabel metal1 1214 1245 1214 1245 1 A_greater_B_node_1
rlabel metal1 1126 1261 1126 1261 1 A3_and_B3c
rlabel metal1 1211 1277 1211 1277 1 A3_nand_B3c
rlabel ndiffusion 1070 1253 1070 1253 1 A_greater_B_node_2
rlabel ndiffusion 1054 1253 1054 1253 1 A_greater_B_node_3
rlabel metal1 1024 1261 1024 1261 1 A3_eq_B3_A2_gt_B2_c
rlabel metal1 969 1279 969 1279 1 A3_eq_B3_A2_gt_B2
rlabel ndiffusion 928 1254 928 1254 1 A_greater_B_node_5
rlabel ndiffusion 907 1255 907 1255 1 A_greater_B_node_6
rlabel ndiffusion 891 1253 891 1253 1 A_greater_B_node_7
rlabel metal1 866 1267 866 1267 1 A3_eq_B3_A2_eq_B2_A1_gt_B1_c
rlabel metal1 812 1280 812 1280 1 A3_eq_B3_A2_eq_B2_A1_gt_B1
rlabel ndiffusion 734 1256 734 1256 1 A_greater_B_node_9
rlabel ndiffusion 715 1255 715 1255 1 A_greater_B_node_10
rlabel ndiffusion 699 1255 699 1255 1 A_greater_B_node_11
rlabel metal1 675 1265 675 1265 1 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c
rlabel metal1 622 1279 622 1279 1 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0
rlabel ndiffusion 750 1254 750 1254 1 A_greater_B_node_8
rlabel pdiffusion 710 1492 710 1492 1 A_GT_B_node_1
rlabel pdiffusion 694 1491 694 1491 1 A_GT_B_node_2
rlabel pdiffusion 677 1493 677 1493 1 A_GT_B_node_3
rlabel metal1 750 1466 750 1466 1 A_GT_B_c
rlabel metal1 792 1483 792 1483 1 A_GT_B
rlabel metal1 948 1547 948 1547 1 A_LS_B_node_1
rlabel metal1 954 1578 954 1578 1 A_LS_B_nand
rlabel metal1 864 1564 864 1564 1 A_LS_B
<< end >>
