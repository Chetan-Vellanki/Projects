magic
tech scmos
timestamp 1701390411
<< nwell >>
rect 863 1035 909 1054
rect 923 1051 984 1068
rect 647 972 731 973
rect 647 953 798 972
rect 809 954 855 973
rect 647 943 752 953
rect 666 769 776 770
rect 855 769 954 770
rect 620 750 776 769
rect 809 750 954 769
rect 967 750 1013 769
rect 674 741 776 750
rect 855 741 954 750
rect 1020 737 1097 769
rect 297 733 361 734
rect 186 714 232 733
rect 257 714 361 733
rect 1125 732 1171 751
rect 1185 748 1246 765
rect 1853 722 1913 739
rect 308 707 361 714
rect 309 706 361 707
rect 1927 706 1973 725
rect 1988 722 2049 739
rect 2063 706 2109 725
rect 2134 724 2195 741
rect 2209 708 2255 727
rect 2282 724 2342 741
rect 2356 708 2402 727
rect 2493 723 2554 740
rect 2568 707 2614 726
rect 2629 723 2690 740
rect 2704 707 2750 726
rect 2775 725 2836 742
rect 2850 709 2896 728
rect 2922 725 2983 742
rect 2997 709 3043 728
rect 376 667 443 695
rect 458 671 504 690
rect 1852 614 1913 631
rect 1927 598 1973 617
rect 1996 614 2057 631
rect 2071 598 2117 617
rect 2145 616 2206 633
rect 2220 600 2266 619
rect 2290 617 2351 634
rect 2365 601 2411 620
rect 1545 544 1606 561
rect 1618 529 1664 548
rect 294 511 358 512
rect 183 492 229 511
rect 254 492 358 511
rect 305 485 358 492
rect 678 486 724 505
rect 738 502 799 519
rect 825 486 871 505
rect 885 502 946 519
rect 306 484 358 485
rect 971 484 1017 503
rect 1031 500 1092 517
rect 1107 484 1153 503
rect 1167 500 1228 517
rect 380 473 403 478
rect 373 445 440 473
rect 455 449 501 468
rect 1544 426 1605 443
rect 669 379 715 398
rect 729 395 790 412
rect 814 378 860 397
rect 874 394 935 411
rect 1617 410 1663 429
rect 963 376 1009 395
rect 1023 392 1084 409
rect 1107 376 1153 395
rect 1167 392 1228 409
rect 1390 390 1474 409
rect 49 338 147 339
rect 3 319 147 338
rect 297 326 361 327
rect 49 310 147 319
rect 161 307 232 326
rect 257 307 361 326
rect 1543 322 1604 339
rect 308 300 361 307
rect 1618 306 1664 325
rect 309 299 361 300
rect 388 291 406 293
rect 383 288 406 291
rect 376 260 443 288
rect 458 264 504 283
rect 1543 226 1604 243
rect 1616 210 1663 229
rect 297 151 361 152
rect 186 132 232 151
rect 257 132 361 151
rect 308 125 361 132
rect 309 124 361 125
rect 379 113 406 118
rect 376 85 443 113
rect 458 89 504 108
<< ntransistor >>
rect 936 1028 941 1033
rect 959 1028 964 1033
rect 878 1020 883 1025
rect 778 938 783 943
rect 835 939 840 944
rect 669 920 674 925
rect 685 920 690 925
rect 701 920 706 925
rect 717 920 722 925
rect 635 735 640 740
rect 824 735 829 740
rect 982 735 987 740
rect 406 717 411 722
rect 424 717 429 722
rect 690 719 695 724
rect 706 719 711 724
rect 722 719 727 724
rect 738 719 743 724
rect 754 719 759 724
rect 883 719 888 724
rect 899 719 904 724
rect 915 719 920 724
rect 931 719 936 724
rect 212 699 217 704
rect 272 699 277 704
rect 1045 718 1050 723
rect 1061 718 1066 723
rect 1077 718 1082 723
rect 1198 725 1203 730
rect 1221 725 1226 730
rect 1140 717 1145 722
rect 1872 699 1877 704
rect 1895 699 1900 704
rect 323 678 328 683
rect 341 678 346 683
rect 2008 699 2013 704
rect 2031 699 2036 704
rect 2154 701 2159 706
rect 2177 701 2182 706
rect 1953 691 1958 696
rect 2089 691 2094 696
rect 2301 701 2306 706
rect 2324 701 2329 706
rect 2235 693 2240 698
rect 2513 700 2518 705
rect 2536 700 2541 705
rect 2382 693 2387 698
rect 2649 700 2654 705
rect 2672 700 2677 705
rect 2795 702 2800 707
rect 2818 702 2823 707
rect 2594 692 2599 697
rect 2730 692 2735 697
rect 2942 702 2947 707
rect 2965 702 2970 707
rect 2876 694 2881 699
rect 3023 694 3028 699
rect 484 656 489 661
rect 1872 591 1877 596
rect 1895 591 1900 596
rect 2016 591 2021 596
rect 2039 591 2044 596
rect 2165 593 2170 598
rect 2188 593 2193 598
rect 2310 594 2315 599
rect 2333 594 2338 599
rect 1953 583 1958 588
rect 2097 583 2102 588
rect 2246 585 2251 590
rect 2391 586 2396 591
rect 1565 521 1570 526
rect 1588 521 1593 526
rect 403 495 408 500
rect 421 495 426 500
rect 209 477 214 482
rect 269 477 274 482
rect 320 456 325 461
rect 338 456 343 461
rect 751 479 756 484
rect 774 479 779 484
rect 693 471 698 476
rect 898 479 903 484
rect 921 479 926 484
rect 1644 514 1649 519
rect 840 471 845 476
rect 1044 477 1049 482
rect 1067 477 1072 482
rect 986 469 991 474
rect 1180 477 1185 482
rect 1203 477 1208 482
rect 1122 469 1127 474
rect 481 434 486 439
rect 742 372 747 377
rect 765 372 770 377
rect 1564 403 1569 408
rect 1587 403 1592 408
rect 684 364 689 369
rect 887 371 892 376
rect 910 371 915 376
rect 1416 375 1421 380
rect 1454 375 1459 380
rect 1643 395 1648 400
rect 829 363 834 368
rect 1036 369 1041 374
rect 1059 369 1064 374
rect 978 361 983 366
rect 1180 369 1185 374
rect 1203 369 1208 374
rect 1122 361 1127 366
rect 18 304 23 309
rect 406 310 411 315
rect 424 310 429 315
rect 1563 299 1568 304
rect 1586 299 1591 304
rect 77 288 82 293
rect 93 288 98 293
rect 109 288 114 293
rect 125 288 130 293
rect 212 292 217 297
rect 272 292 277 297
rect 323 271 328 276
rect 341 271 346 276
rect 1644 291 1649 296
rect 484 249 489 254
rect 1563 203 1568 208
rect 1586 203 1591 208
rect 1643 195 1648 200
rect 406 135 411 140
rect 424 135 429 140
rect 212 117 217 122
rect 272 117 277 122
rect 323 96 328 101
rect 341 96 346 101
rect 484 74 489 79
<< ptransistor >>
rect 936 1057 941 1062
rect 959 1057 964 1062
rect 878 1042 883 1047
rect 669 956 674 961
rect 685 956 690 961
rect 701 956 706 961
rect 717 956 722 961
rect 778 960 783 965
rect 835 961 840 966
rect 635 757 640 762
rect 690 753 695 758
rect 706 753 711 758
rect 722 753 727 758
rect 738 753 743 758
rect 754 753 759 758
rect 824 757 829 762
rect 212 721 217 726
rect 272 721 277 726
rect 883 753 888 758
rect 899 753 904 758
rect 915 753 920 758
rect 931 753 936 758
rect 982 757 987 762
rect 1045 752 1050 757
rect 1061 752 1066 757
rect 1077 752 1082 757
rect 1198 754 1203 759
rect 1221 754 1226 759
rect 323 717 328 722
rect 341 717 346 722
rect 1140 739 1145 744
rect 1872 728 1877 733
rect 1895 728 1900 733
rect 2008 728 2013 733
rect 2031 728 2036 733
rect 2154 730 2159 735
rect 2177 730 2182 735
rect 2301 730 2306 735
rect 2324 730 2329 735
rect 1953 713 1958 718
rect 2089 713 2094 718
rect 2235 715 2240 720
rect 2513 729 2518 734
rect 2536 729 2541 734
rect 2649 729 2654 734
rect 2672 729 2677 734
rect 2795 731 2800 736
rect 2818 731 2823 736
rect 2942 731 2947 736
rect 2965 731 2970 736
rect 2382 715 2387 720
rect 406 678 411 683
rect 424 678 429 683
rect 484 678 489 683
rect 2594 714 2599 719
rect 2730 714 2735 719
rect 2876 716 2881 721
rect 3023 716 3028 721
rect 1872 620 1877 625
rect 1895 620 1900 625
rect 2016 620 2021 625
rect 2039 620 2044 625
rect 2165 622 2170 627
rect 2188 622 2193 627
rect 2310 623 2315 628
rect 2333 623 2338 628
rect 1953 605 1958 610
rect 2097 605 2102 610
rect 2246 607 2251 612
rect 2391 608 2396 613
rect 1565 550 1570 555
rect 1588 550 1593 555
rect 209 499 214 504
rect 269 499 274 504
rect 1644 536 1649 541
rect 751 508 756 513
rect 774 508 779 513
rect 898 508 903 513
rect 921 508 926 513
rect 320 495 325 500
rect 338 495 343 500
rect 693 493 698 498
rect 840 493 845 498
rect 1044 506 1049 511
rect 1067 506 1072 511
rect 1180 506 1185 511
rect 1203 506 1208 511
rect 986 491 991 496
rect 403 456 408 461
rect 421 456 426 461
rect 481 456 486 461
rect 1122 491 1127 496
rect 1564 432 1569 437
rect 1587 432 1592 437
rect 742 401 747 406
rect 765 401 770 406
rect 684 386 689 391
rect 887 400 892 405
rect 910 400 915 405
rect 1643 417 1648 422
rect 829 385 834 390
rect 1036 398 1041 403
rect 1059 398 1064 403
rect 1180 398 1185 403
rect 1203 398 1208 403
rect 978 383 983 388
rect 1122 383 1127 388
rect 1416 397 1421 402
rect 1454 397 1459 402
rect 18 326 23 331
rect 77 322 82 327
rect 93 322 98 327
rect 109 322 114 327
rect 125 322 130 327
rect 212 314 217 319
rect 272 314 277 319
rect 1563 328 1568 333
rect 1586 328 1591 333
rect 323 310 328 315
rect 341 310 346 315
rect 1644 313 1649 318
rect 406 271 411 276
rect 424 271 429 276
rect 484 271 489 276
rect 1563 232 1568 237
rect 1586 232 1591 237
rect 1643 217 1648 222
rect 212 139 217 144
rect 272 139 277 144
rect 323 135 328 140
rect 341 135 346 140
rect 406 96 411 101
rect 424 96 429 101
rect 484 96 489 101
<< ndiffusion >>
rect 934 1028 936 1033
rect 941 1028 943 1033
rect 957 1028 959 1033
rect 964 1028 966 1033
rect 875 1020 878 1025
rect 883 1020 885 1025
rect 776 938 778 943
rect 783 938 786 943
rect 833 939 835 944
rect 840 939 843 944
rect 666 920 669 925
rect 674 920 677 925
rect 682 920 685 925
rect 690 920 693 925
rect 698 920 701 925
rect 706 920 709 925
rect 714 920 717 925
rect 722 920 725 925
rect 632 735 635 740
rect 640 735 642 740
rect 821 735 824 740
rect 829 735 831 740
rect 979 735 982 740
rect 987 735 989 740
rect 403 717 406 722
rect 411 717 424 722
rect 429 717 432 722
rect 687 719 690 724
rect 695 719 706 724
rect 711 719 722 724
rect 727 719 738 724
rect 743 719 754 724
rect 759 719 762 724
rect 881 719 883 724
rect 888 719 899 724
rect 904 719 915 724
rect 920 719 931 724
rect 936 719 939 724
rect 210 699 212 704
rect 217 699 220 704
rect 269 699 272 704
rect 277 699 279 704
rect 1039 718 1045 723
rect 1050 718 1061 723
rect 1066 718 1077 723
rect 1082 718 1085 723
rect 1196 725 1198 730
rect 1203 725 1205 730
rect 1219 725 1221 730
rect 1226 725 1228 730
rect 1137 717 1140 722
rect 1145 717 1147 722
rect 1870 699 1872 704
rect 1877 699 1879 704
rect 1893 699 1895 704
rect 1900 699 1902 704
rect 320 678 323 683
rect 328 678 341 683
rect 346 678 349 683
rect 2006 699 2008 704
rect 2013 699 2015 704
rect 2029 699 2031 704
rect 2036 699 2038 704
rect 2152 701 2154 706
rect 2159 701 2161 706
rect 2175 701 2177 706
rect 2182 701 2184 706
rect 1951 691 1953 696
rect 1958 691 1961 696
rect 2087 691 2089 696
rect 2094 691 2097 696
rect 2299 701 2301 706
rect 2306 701 2308 706
rect 2322 701 2324 706
rect 2329 701 2331 706
rect 2233 693 2235 698
rect 2240 693 2243 698
rect 2511 700 2513 705
rect 2518 700 2520 705
rect 2534 700 2536 705
rect 2541 700 2543 705
rect 2380 693 2382 698
rect 2387 693 2390 698
rect 2647 700 2649 705
rect 2654 700 2656 705
rect 2670 700 2672 705
rect 2677 700 2679 705
rect 2793 702 2795 707
rect 2800 702 2802 707
rect 2816 702 2818 707
rect 2823 702 2825 707
rect 2592 692 2594 697
rect 2599 692 2602 697
rect 2728 692 2730 697
rect 2735 692 2738 697
rect 2940 702 2942 707
rect 2947 702 2949 707
rect 2963 702 2965 707
rect 2970 702 2972 707
rect 2874 694 2876 699
rect 2881 694 2884 699
rect 3021 694 3023 699
rect 3028 694 3031 699
rect 482 656 484 661
rect 489 656 492 661
rect 1870 591 1872 596
rect 1877 591 1879 596
rect 1893 591 1895 596
rect 1900 591 1902 596
rect 2014 591 2016 596
rect 2021 591 2023 596
rect 2037 591 2039 596
rect 2044 591 2046 596
rect 2163 593 2165 598
rect 2170 593 2172 598
rect 2186 593 2188 598
rect 2193 593 2195 598
rect 2308 594 2310 599
rect 2315 594 2317 599
rect 2331 594 2333 599
rect 2338 594 2340 599
rect 1951 583 1953 588
rect 1958 583 1961 588
rect 2095 583 2097 588
rect 2102 583 2105 588
rect 2244 585 2246 590
rect 2251 585 2254 590
rect 2389 586 2391 591
rect 2396 586 2399 591
rect 1563 521 1565 526
rect 1570 521 1572 526
rect 1586 521 1588 526
rect 1593 521 1595 526
rect 400 495 403 500
rect 408 495 421 500
rect 426 495 429 500
rect 207 477 209 482
rect 214 477 217 482
rect 266 477 269 482
rect 274 477 276 482
rect 317 456 320 461
rect 325 456 338 461
rect 343 456 346 461
rect 749 479 751 484
rect 756 479 758 484
rect 772 479 774 484
rect 779 479 781 484
rect 690 471 693 476
rect 698 471 700 476
rect 896 479 898 484
rect 903 479 905 484
rect 919 479 921 484
rect 926 479 928 484
rect 1642 514 1644 519
rect 1649 514 1652 519
rect 837 471 840 476
rect 845 471 847 476
rect 1042 477 1044 482
rect 1049 477 1051 482
rect 1065 477 1067 482
rect 1072 477 1074 482
rect 983 469 986 474
rect 991 469 993 474
rect 1178 477 1180 482
rect 1185 477 1187 482
rect 1201 477 1203 482
rect 1208 477 1210 482
rect 1119 469 1122 474
rect 1127 469 1129 474
rect 479 434 481 439
rect 486 434 489 439
rect 740 372 742 377
rect 747 372 749 377
rect 763 372 765 377
rect 770 372 772 377
rect 1562 403 1564 408
rect 1569 403 1571 408
rect 1585 403 1587 408
rect 1592 403 1594 408
rect 681 364 684 369
rect 689 364 691 369
rect 885 371 887 376
rect 892 371 894 376
rect 908 371 910 376
rect 915 371 917 376
rect 1414 375 1416 380
rect 1421 375 1424 380
rect 1452 375 1454 380
rect 1459 375 1462 380
rect 1641 395 1643 400
rect 1648 395 1651 400
rect 826 363 829 368
rect 834 363 836 368
rect 1034 369 1036 374
rect 1041 369 1043 374
rect 1057 369 1059 374
rect 1064 369 1066 374
rect 975 361 978 366
rect 983 361 985 366
rect 1178 369 1180 374
rect 1185 369 1187 374
rect 1201 369 1203 374
rect 1208 369 1210 374
rect 1119 361 1122 366
rect 1127 361 1129 366
rect 15 304 18 309
rect 23 304 25 309
rect 403 310 406 315
rect 411 310 424 315
rect 429 310 432 315
rect 1561 299 1563 304
rect 1568 299 1570 304
rect 1584 299 1586 304
rect 1591 299 1593 304
rect 75 288 77 293
rect 82 288 93 293
rect 98 288 109 293
rect 114 288 125 293
rect 130 288 133 293
rect 210 292 212 297
rect 217 292 220 297
rect 269 292 272 297
rect 277 292 279 297
rect 320 271 323 276
rect 328 271 341 276
rect 346 271 349 276
rect 1642 291 1644 296
rect 1649 291 1652 296
rect 482 249 484 254
rect 489 249 492 254
rect 1561 203 1563 208
rect 1568 203 1570 208
rect 1584 203 1586 208
rect 1591 203 1593 208
rect 1641 195 1643 200
rect 1648 195 1651 200
rect 403 135 406 140
rect 411 135 424 140
rect 429 135 432 140
rect 210 117 212 122
rect 217 117 220 122
rect 269 117 272 122
rect 277 117 279 122
rect 320 96 323 101
rect 328 96 341 101
rect 346 96 349 101
rect 482 74 484 79
rect 489 74 492 79
<< pdiffusion >>
rect 934 1057 936 1062
rect 941 1057 947 1062
rect 952 1057 959 1062
rect 964 1057 966 1062
rect 875 1042 878 1047
rect 883 1042 885 1047
rect 666 956 669 961
rect 674 956 685 961
rect 690 956 701 961
rect 706 956 717 961
rect 722 956 725 961
rect 776 960 778 965
rect 783 960 786 965
rect 833 961 835 966
rect 840 961 843 966
rect 632 757 635 762
rect 640 757 642 762
rect 687 753 690 758
rect 695 753 698 758
rect 703 753 706 758
rect 711 753 714 758
rect 719 753 722 758
rect 727 753 730 758
rect 735 753 738 758
rect 743 753 746 758
rect 751 753 754 758
rect 759 753 762 758
rect 821 757 824 762
rect 829 757 831 762
rect 210 721 212 726
rect 217 721 220 726
rect 269 721 272 726
rect 277 721 279 726
rect 880 753 883 758
rect 888 753 891 758
rect 896 753 899 758
rect 904 753 907 758
rect 912 753 915 758
rect 920 753 923 758
rect 928 753 931 758
rect 936 753 939 758
rect 979 757 982 762
rect 987 757 989 762
rect 1042 752 1045 757
rect 1050 752 1053 757
rect 1058 752 1061 757
rect 1066 752 1069 757
rect 1074 752 1077 757
rect 1082 752 1085 757
rect 1196 754 1198 759
rect 1203 754 1209 759
rect 1214 754 1221 759
rect 1226 754 1228 759
rect 320 717 323 722
rect 328 717 341 722
rect 346 717 349 722
rect 1137 739 1140 744
rect 1145 739 1147 744
rect 1870 728 1872 733
rect 1877 728 1884 733
rect 1889 728 1895 733
rect 1900 728 1902 733
rect 2006 728 2008 733
rect 2013 728 2020 733
rect 2025 728 2031 733
rect 2036 728 2038 733
rect 2152 730 2154 735
rect 2159 730 2166 735
rect 2171 730 2177 735
rect 2182 730 2184 735
rect 2299 730 2301 735
rect 2306 730 2313 735
rect 2318 730 2324 735
rect 2329 730 2331 735
rect 1951 713 1953 718
rect 1958 713 1961 718
rect 2087 713 2089 718
rect 2094 713 2097 718
rect 2233 715 2235 720
rect 2240 715 2243 720
rect 2511 729 2513 734
rect 2518 729 2525 734
rect 2530 729 2536 734
rect 2541 729 2543 734
rect 2647 729 2649 734
rect 2654 729 2661 734
rect 2666 729 2672 734
rect 2677 729 2679 734
rect 2793 731 2795 736
rect 2800 731 2807 736
rect 2812 731 2818 736
rect 2823 731 2825 736
rect 2940 731 2942 736
rect 2947 731 2954 736
rect 2959 731 2965 736
rect 2970 731 2972 736
rect 2380 715 2382 720
rect 2387 715 2390 720
rect 403 678 406 683
rect 411 678 424 683
rect 429 678 432 683
rect 482 678 484 683
rect 489 678 492 683
rect 2592 714 2594 719
rect 2599 714 2602 719
rect 2728 714 2730 719
rect 2735 714 2738 719
rect 2874 716 2876 721
rect 2881 716 2884 721
rect 3021 716 3023 721
rect 3028 716 3031 721
rect 1870 620 1872 625
rect 1877 620 1884 625
rect 1889 620 1895 625
rect 1900 620 1902 625
rect 2014 620 2016 625
rect 2021 620 2028 625
rect 2033 620 2039 625
rect 2044 620 2046 625
rect 2163 622 2165 627
rect 2170 622 2177 627
rect 2182 622 2188 627
rect 2193 622 2195 627
rect 2308 623 2310 628
rect 2315 623 2322 628
rect 2327 623 2333 628
rect 2338 623 2340 628
rect 1951 605 1953 610
rect 1958 605 1961 610
rect 2095 605 2097 610
rect 2102 605 2105 610
rect 2244 607 2246 612
rect 2251 607 2254 612
rect 2389 608 2391 613
rect 2396 608 2399 613
rect 1563 550 1565 555
rect 1570 550 1577 555
rect 1582 550 1588 555
rect 1593 550 1595 555
rect 207 499 209 504
rect 214 499 217 504
rect 266 499 269 504
rect 274 499 276 504
rect 1642 536 1644 541
rect 1649 536 1652 541
rect 749 508 751 513
rect 756 508 762 513
rect 767 508 774 513
rect 779 508 781 513
rect 896 508 898 513
rect 903 508 909 513
rect 914 508 921 513
rect 926 508 928 513
rect 317 495 320 500
rect 325 495 338 500
rect 343 495 346 500
rect 690 493 693 498
rect 698 493 700 498
rect 837 493 840 498
rect 845 493 847 498
rect 1042 506 1044 511
rect 1049 506 1055 511
rect 1060 506 1067 511
rect 1072 506 1074 511
rect 1178 506 1180 511
rect 1185 506 1191 511
rect 1196 506 1203 511
rect 1208 506 1210 511
rect 983 491 986 496
rect 991 491 993 496
rect 400 456 403 461
rect 408 456 421 461
rect 426 456 429 461
rect 479 456 481 461
rect 486 456 489 461
rect 1119 491 1122 496
rect 1127 491 1129 496
rect 1562 432 1564 437
rect 1569 432 1576 437
rect 1581 432 1587 437
rect 1592 432 1594 437
rect 740 401 742 406
rect 747 401 753 406
rect 758 401 765 406
rect 770 401 772 406
rect 681 386 684 391
rect 689 386 691 391
rect 885 400 887 405
rect 892 400 898 405
rect 903 400 910 405
rect 915 400 917 405
rect 1641 417 1643 422
rect 1648 417 1651 422
rect 826 385 829 390
rect 834 385 836 390
rect 1034 398 1036 403
rect 1041 398 1047 403
rect 1052 398 1059 403
rect 1064 398 1066 403
rect 1178 398 1180 403
rect 1185 398 1191 403
rect 1196 398 1203 403
rect 1208 398 1210 403
rect 975 383 978 388
rect 983 383 985 388
rect 1119 383 1122 388
rect 1127 383 1129 388
rect 1414 397 1416 402
rect 1421 397 1424 402
rect 1452 397 1454 402
rect 1459 397 1462 402
rect 15 326 18 331
rect 23 326 25 331
rect 74 322 77 327
rect 82 322 85 327
rect 90 322 93 327
rect 98 322 101 327
rect 106 322 109 327
rect 114 322 117 327
rect 122 322 125 327
rect 130 322 133 327
rect 210 314 212 319
rect 217 314 220 319
rect 269 314 272 319
rect 277 314 279 319
rect 1561 328 1563 333
rect 1568 328 1575 333
rect 1580 328 1586 333
rect 1591 328 1593 333
rect 320 310 323 315
rect 328 310 341 315
rect 346 310 349 315
rect 1642 313 1644 318
rect 1649 313 1652 318
rect 403 271 406 276
rect 411 271 424 276
rect 429 271 432 276
rect 482 271 484 276
rect 489 271 492 276
rect 1561 232 1563 237
rect 1568 232 1575 237
rect 1580 232 1586 237
rect 1591 232 1593 237
rect 1641 217 1643 222
rect 1648 217 1651 222
rect 210 139 212 144
rect 217 139 220 144
rect 269 139 272 144
rect 277 139 279 144
rect 320 135 323 140
rect 328 135 341 140
rect 346 135 349 140
rect 403 96 406 101
rect 411 96 424 101
rect 429 96 432 101
rect 482 96 484 101
rect 489 96 492 101
<< ndcontact >>
rect 929 1028 934 1033
rect 943 1028 947 1033
rect 953 1028 957 1033
rect 966 1028 971 1033
rect 870 1020 875 1025
rect 885 1020 890 1025
rect 771 938 776 943
rect 786 938 791 943
rect 828 939 833 944
rect 843 939 848 944
rect 661 920 666 925
rect 677 920 682 925
rect 693 920 698 925
rect 709 920 714 925
rect 725 920 730 925
rect 627 735 632 740
rect 642 735 647 740
rect 816 735 821 740
rect 831 735 836 740
rect 974 735 979 740
rect 989 735 994 740
rect 398 717 403 722
rect 432 717 437 722
rect 682 719 687 724
rect 762 719 767 724
rect 876 719 881 724
rect 939 719 944 724
rect 205 699 210 704
rect 220 699 225 704
rect 264 699 269 704
rect 279 699 284 704
rect 1034 718 1039 723
rect 1085 718 1090 723
rect 1191 725 1196 730
rect 1205 725 1209 730
rect 1215 725 1219 730
rect 1228 725 1233 730
rect 1132 717 1137 722
rect 1147 717 1152 722
rect 1865 699 1870 704
rect 1879 699 1883 704
rect 1889 699 1893 704
rect 1902 699 1907 704
rect 315 678 320 683
rect 349 678 354 683
rect 2001 699 2006 704
rect 2015 699 2019 704
rect 2025 699 2029 704
rect 2038 699 2043 704
rect 2147 701 2152 706
rect 2161 701 2165 706
rect 2171 701 2175 706
rect 2184 701 2189 706
rect 1946 691 1951 696
rect 1961 691 1966 696
rect 2082 691 2087 696
rect 2097 691 2102 696
rect 2294 701 2299 706
rect 2308 701 2312 706
rect 2318 701 2322 706
rect 2331 701 2336 706
rect 2228 693 2233 698
rect 2243 693 2248 698
rect 2506 700 2511 705
rect 2520 700 2524 705
rect 2530 700 2534 705
rect 2543 700 2548 705
rect 2375 693 2380 698
rect 2390 693 2395 698
rect 2642 700 2647 705
rect 2656 700 2660 705
rect 2666 700 2670 705
rect 2679 700 2684 705
rect 2788 702 2793 707
rect 2802 702 2806 707
rect 2812 702 2816 707
rect 2825 702 2830 707
rect 2587 692 2592 697
rect 2602 692 2607 697
rect 2723 692 2728 697
rect 2738 692 2743 697
rect 2935 702 2940 707
rect 2949 702 2953 707
rect 2959 702 2963 707
rect 2972 702 2977 707
rect 2869 694 2874 699
rect 2884 694 2889 699
rect 3016 694 3021 699
rect 3031 694 3036 699
rect 477 656 482 661
rect 492 656 497 661
rect 1865 591 1870 596
rect 1879 591 1883 596
rect 1889 591 1893 596
rect 1902 591 1907 596
rect 2009 591 2014 596
rect 2023 591 2027 596
rect 2033 591 2037 596
rect 2046 591 2051 596
rect 2158 593 2163 598
rect 2172 593 2176 598
rect 2182 593 2186 598
rect 2195 593 2200 598
rect 2303 594 2308 599
rect 2317 594 2321 599
rect 2327 594 2331 599
rect 2340 594 2345 599
rect 1946 583 1951 588
rect 1961 583 1966 588
rect 2090 583 2095 588
rect 2105 583 2110 588
rect 2239 585 2244 590
rect 2254 585 2259 590
rect 2384 586 2389 591
rect 2399 586 2404 591
rect 1558 521 1563 526
rect 1572 521 1576 526
rect 1582 521 1586 526
rect 1595 521 1600 526
rect 395 495 400 500
rect 429 495 434 500
rect 202 477 207 482
rect 217 477 222 482
rect 261 477 266 482
rect 276 477 281 482
rect 312 456 317 461
rect 346 456 351 461
rect 744 479 749 484
rect 758 479 762 484
rect 768 479 772 484
rect 781 479 786 484
rect 685 471 690 476
rect 700 471 705 476
rect 891 479 896 484
rect 905 479 909 484
rect 915 479 919 484
rect 928 479 933 484
rect 1637 514 1642 519
rect 1652 514 1657 519
rect 832 471 837 476
rect 847 471 852 476
rect 1037 477 1042 482
rect 1051 477 1055 482
rect 1061 477 1065 482
rect 1074 477 1079 482
rect 978 469 983 474
rect 993 469 998 474
rect 1173 477 1178 482
rect 1187 477 1191 482
rect 1197 477 1201 482
rect 1210 477 1215 482
rect 1114 469 1119 474
rect 1129 469 1134 474
rect 474 434 479 439
rect 489 434 494 439
rect 735 372 740 377
rect 749 372 753 377
rect 759 372 763 377
rect 772 372 777 377
rect 1557 403 1562 408
rect 1571 403 1575 408
rect 1581 403 1585 408
rect 1594 403 1599 408
rect 676 364 681 369
rect 691 364 696 369
rect 880 371 885 376
rect 894 371 898 376
rect 904 371 908 376
rect 917 371 922 376
rect 1409 375 1414 380
rect 1424 375 1429 380
rect 1447 375 1452 380
rect 1462 375 1467 380
rect 1636 395 1641 400
rect 1651 395 1656 400
rect 821 363 826 368
rect 836 363 841 368
rect 1029 369 1034 374
rect 1043 369 1047 374
rect 1053 369 1057 374
rect 1066 369 1071 374
rect 970 361 975 366
rect 985 361 990 366
rect 1173 369 1178 374
rect 1187 369 1191 374
rect 1197 369 1201 374
rect 1210 369 1215 374
rect 1114 361 1119 366
rect 1129 361 1134 366
rect 10 304 15 309
rect 25 304 30 309
rect 398 310 403 315
rect 432 310 437 315
rect 1556 299 1561 304
rect 1570 299 1574 304
rect 1580 299 1584 304
rect 1593 299 1598 304
rect 70 288 75 293
rect 133 288 138 293
rect 205 292 210 297
rect 220 292 225 297
rect 264 292 269 297
rect 279 292 284 297
rect 315 271 320 276
rect 349 271 354 276
rect 1637 291 1642 296
rect 1652 291 1657 296
rect 477 249 482 254
rect 492 249 497 254
rect 1556 203 1561 208
rect 1570 203 1574 208
rect 1580 203 1584 208
rect 1593 203 1598 208
rect 1636 195 1641 200
rect 1651 195 1656 200
rect 398 135 403 140
rect 432 135 437 140
rect 205 117 210 122
rect 220 117 225 122
rect 264 117 269 122
rect 279 117 284 122
rect 315 96 320 101
rect 349 96 354 101
rect 477 74 482 79
rect 492 74 497 79
<< pdcontact >>
rect 929 1057 934 1062
rect 947 1057 952 1062
rect 966 1057 971 1062
rect 870 1042 875 1047
rect 885 1042 890 1047
rect 661 956 666 961
rect 725 956 730 961
rect 771 960 776 965
rect 786 960 791 965
rect 828 961 833 966
rect 843 961 848 966
rect 627 757 632 762
rect 642 757 647 762
rect 682 753 687 758
rect 698 753 703 758
rect 714 753 719 758
rect 730 753 735 758
rect 746 753 751 758
rect 762 753 767 758
rect 816 757 821 762
rect 831 757 836 762
rect 205 721 210 726
rect 220 721 225 726
rect 264 721 269 726
rect 279 721 284 726
rect 875 753 880 758
rect 891 753 896 758
rect 907 753 912 758
rect 923 753 928 758
rect 939 753 944 758
rect 974 757 979 762
rect 989 757 994 762
rect 1037 752 1042 757
rect 1053 752 1058 757
rect 1069 752 1074 757
rect 1085 752 1090 757
rect 1191 754 1196 759
rect 1209 754 1214 759
rect 1228 754 1233 759
rect 315 717 320 722
rect 349 717 354 722
rect 1132 739 1137 744
rect 1147 739 1152 744
rect 1865 728 1870 733
rect 1884 728 1889 733
rect 1902 728 1907 733
rect 2001 728 2006 733
rect 2020 728 2025 733
rect 2038 728 2043 733
rect 2147 730 2152 735
rect 2166 730 2171 735
rect 2184 730 2189 735
rect 2294 730 2299 735
rect 2313 730 2318 735
rect 2331 730 2336 735
rect 1946 713 1951 718
rect 1961 713 1966 718
rect 2082 713 2087 718
rect 2097 713 2102 718
rect 2228 715 2233 720
rect 2243 715 2248 720
rect 2506 729 2511 734
rect 2525 729 2530 734
rect 2543 729 2548 734
rect 2642 729 2647 734
rect 2661 729 2666 734
rect 2679 729 2684 734
rect 2788 731 2793 736
rect 2807 731 2812 736
rect 2825 731 2830 736
rect 2935 731 2940 736
rect 2954 731 2959 736
rect 2972 731 2977 736
rect 2375 715 2380 720
rect 2390 715 2395 720
rect 398 678 403 683
rect 432 678 437 683
rect 477 678 482 683
rect 492 678 497 683
rect 2587 714 2592 719
rect 2602 714 2607 719
rect 2723 714 2728 719
rect 2738 714 2743 719
rect 2869 716 2874 721
rect 2884 716 2889 721
rect 3016 716 3021 721
rect 3031 716 3036 721
rect 1865 620 1870 625
rect 1884 620 1889 625
rect 1902 620 1907 625
rect 2009 620 2014 625
rect 2028 620 2033 625
rect 2046 620 2051 625
rect 2158 622 2163 627
rect 2177 622 2182 627
rect 2195 622 2200 627
rect 2303 623 2308 628
rect 2322 623 2327 628
rect 2340 623 2345 628
rect 1946 605 1951 610
rect 1961 605 1966 610
rect 2090 605 2095 610
rect 2105 605 2110 610
rect 2239 607 2244 612
rect 2254 607 2259 612
rect 2384 608 2389 613
rect 2399 608 2404 613
rect 1558 550 1563 555
rect 1577 550 1582 555
rect 1595 550 1600 555
rect 202 499 207 504
rect 217 499 222 504
rect 261 499 266 504
rect 276 499 281 504
rect 1637 536 1642 541
rect 1652 536 1657 541
rect 744 508 749 513
rect 762 508 767 513
rect 781 508 786 513
rect 891 508 896 513
rect 909 508 914 513
rect 928 508 933 513
rect 312 495 317 500
rect 346 495 351 500
rect 685 493 690 498
rect 700 493 705 498
rect 832 493 837 498
rect 847 493 852 498
rect 1037 506 1042 511
rect 1055 506 1060 511
rect 1074 506 1079 511
rect 1173 506 1178 511
rect 1191 506 1196 511
rect 1210 506 1215 511
rect 978 491 983 496
rect 993 491 998 496
rect 395 456 400 461
rect 429 456 434 461
rect 474 456 479 461
rect 489 456 494 461
rect 1114 491 1119 496
rect 1129 491 1134 496
rect 1557 432 1562 437
rect 1576 432 1581 437
rect 1594 432 1599 437
rect 735 401 740 406
rect 753 401 758 406
rect 772 401 777 406
rect 676 386 681 391
rect 691 386 696 391
rect 880 400 885 405
rect 898 400 903 405
rect 917 400 922 405
rect 1636 417 1641 422
rect 1651 417 1656 422
rect 821 385 826 390
rect 836 385 841 390
rect 1029 398 1034 403
rect 1047 398 1052 403
rect 1066 398 1071 403
rect 1173 398 1178 403
rect 1191 398 1196 403
rect 1210 398 1215 403
rect 970 383 975 388
rect 985 383 990 388
rect 1114 383 1119 388
rect 1129 383 1134 388
rect 1409 397 1414 402
rect 1424 397 1429 402
rect 1447 397 1452 402
rect 1462 397 1467 402
rect 10 326 15 331
rect 25 326 30 331
rect 69 322 74 327
rect 85 322 90 327
rect 101 322 106 327
rect 117 322 122 327
rect 133 322 138 327
rect 205 314 210 319
rect 220 314 225 319
rect 264 314 269 319
rect 279 314 284 319
rect 1556 328 1561 333
rect 1575 328 1580 333
rect 1593 328 1598 333
rect 315 310 320 315
rect 349 310 354 315
rect 1637 313 1642 318
rect 1652 313 1657 318
rect 398 271 403 276
rect 432 271 437 276
rect 477 271 482 276
rect 492 271 497 276
rect 1556 232 1561 237
rect 1575 232 1580 237
rect 1593 232 1598 237
rect 1636 217 1641 222
rect 1651 217 1656 222
rect 205 139 210 144
rect 220 139 225 144
rect 264 139 269 144
rect 279 139 284 144
rect 315 135 320 140
rect 349 135 354 140
rect 398 96 403 101
rect 432 96 437 101
rect 477 96 482 101
rect 492 96 497 101
<< nsubstratencontact >>
rect 975 1057 980 1062
rect 897 1042 902 1047
rect 737 956 742 961
rect 759 960 764 965
rect 816 961 821 966
rect 654 757 659 762
rect 843 757 848 762
rect 193 721 198 726
rect 291 721 296 726
rect 863 753 868 758
rect 1001 757 1006 762
rect 1027 752 1032 757
rect 1237 754 1242 759
rect 303 717 308 722
rect 1159 739 1164 744
rect 1856 728 1861 733
rect 1992 728 1997 733
rect 2139 730 2143 735
rect 2285 730 2290 735
rect 1934 713 1939 718
rect 2070 713 2075 718
rect 2216 715 2221 720
rect 2497 729 2502 734
rect 2633 729 2638 734
rect 2779 731 2784 736
rect 2926 731 2931 736
rect 2363 715 2368 720
rect 383 676 389 682
rect 465 678 470 683
rect 2575 714 2580 719
rect 2711 714 2716 719
rect 2857 716 2862 721
rect 3004 716 3009 721
rect 1856 620 1861 625
rect 2000 620 2005 625
rect 2149 622 2154 627
rect 2294 623 2299 628
rect 1934 605 1939 610
rect 2078 605 2083 610
rect 2227 607 2232 612
rect 2372 608 2377 613
rect 1549 550 1554 555
rect 190 499 195 504
rect 288 499 293 504
rect 1625 536 1630 541
rect 790 508 795 513
rect 937 508 942 513
rect 300 495 305 500
rect 712 493 717 498
rect 859 493 864 498
rect 1083 506 1088 511
rect 1219 506 1224 511
rect 1005 491 1010 496
rect 380 457 386 462
rect 462 456 467 461
rect 1141 491 1146 496
rect 1548 432 1553 437
rect 781 401 786 406
rect 703 386 708 391
rect 926 400 931 405
rect 1624 417 1629 422
rect 848 385 853 390
rect 1075 398 1080 403
rect 1219 398 1224 403
rect 997 383 1002 388
rect 1141 383 1146 388
rect 1397 397 1402 402
rect 37 326 42 331
rect 57 322 62 327
rect 168 314 173 319
rect 291 314 296 319
rect 1547 328 1552 333
rect 303 310 308 315
rect 1625 313 1630 318
rect 383 269 388 275
rect 465 271 470 276
rect 1547 232 1552 237
rect 1624 217 1629 222
rect 193 139 198 144
rect 291 139 296 144
rect 303 135 308 140
rect 383 96 388 101
rect 465 96 470 101
<< polysilicon >>
rect 936 1062 941 1076
rect 959 1062 964 1076
rect 878 1047 883 1050
rect 878 1033 883 1042
rect 936 1033 941 1057
rect 959 1033 964 1057
rect 878 1029 882 1033
rect 878 1025 883 1029
rect 878 1015 883 1020
rect 936 1009 941 1028
rect 959 1009 964 1028
rect 778 965 783 968
rect 835 966 840 969
rect 669 961 674 964
rect 685 961 690 964
rect 701 961 706 964
rect 717 961 722 964
rect 669 925 674 956
rect 685 925 690 956
rect 701 925 706 956
rect 717 925 722 956
rect 778 951 783 960
rect 835 952 840 961
rect 779 947 783 951
rect 836 948 840 952
rect 778 943 783 947
rect 835 944 840 948
rect 778 933 783 938
rect 835 934 840 939
rect 669 909 674 920
rect 685 909 690 920
rect 701 909 706 920
rect 717 910 722 920
rect 635 762 640 765
rect 690 758 695 762
rect 706 758 711 762
rect 722 758 727 777
rect 738 758 743 777
rect 824 762 829 765
rect 754 758 759 762
rect 635 748 640 757
rect 883 758 888 777
rect 899 758 904 777
rect 915 758 920 762
rect 931 758 936 777
rect 982 762 987 765
rect 341 743 379 744
rect 635 744 639 748
rect 384 743 429 744
rect 341 739 429 743
rect 635 740 640 744
rect 212 726 217 729
rect 272 726 277 729
rect 323 722 328 726
rect 341 722 346 739
rect 406 722 411 726
rect 424 722 429 739
rect 635 730 640 735
rect 690 724 695 753
rect 706 724 711 753
rect 722 724 727 753
rect 738 724 743 753
rect 754 724 759 753
rect 824 748 829 757
rect 1045 757 1050 762
rect 1061 757 1066 779
rect 1077 757 1082 777
rect 1198 759 1203 773
rect 1221 759 1226 773
rect 824 744 828 748
rect 824 740 829 744
rect 824 730 829 735
rect 883 724 888 753
rect 899 724 904 753
rect 915 724 920 753
rect 931 724 936 753
rect 982 748 987 757
rect 982 744 986 748
rect 982 740 987 744
rect 982 730 987 735
rect 212 712 217 721
rect 213 708 217 712
rect 212 704 217 708
rect 272 712 277 721
rect 1045 723 1050 752
rect 1061 723 1066 752
rect 1077 723 1082 752
rect 1140 744 1145 747
rect 1140 730 1145 739
rect 1198 730 1203 754
rect 1221 730 1226 754
rect 1872 733 1877 747
rect 1895 733 1900 747
rect 2008 733 2013 747
rect 2031 733 2036 747
rect 2154 735 2159 749
rect 2177 735 2182 749
rect 2301 735 2306 749
rect 2324 735 2329 749
rect 1140 726 1144 730
rect 272 708 276 712
rect 272 704 277 708
rect 323 705 328 717
rect 341 713 346 717
rect 406 705 411 717
rect 424 713 429 717
rect 324 700 346 705
rect 406 700 429 705
rect 690 700 695 719
rect 212 694 217 699
rect 272 694 277 699
rect 304 688 328 693
rect 304 680 309 688
rect 323 683 328 688
rect 341 683 346 700
rect 406 683 411 687
rect 424 683 429 700
rect 706 699 711 719
rect 722 702 727 719
rect 738 702 743 719
rect 754 699 759 719
rect 883 712 888 719
rect 899 712 904 719
rect 915 702 920 719
rect 931 702 936 719
rect 1140 722 1145 726
rect 2513 734 2518 748
rect 2536 734 2541 748
rect 2649 734 2654 748
rect 2672 734 2677 748
rect 2795 736 2800 750
rect 2818 736 2823 750
rect 2942 736 2947 750
rect 2965 736 2970 750
rect 1045 703 1050 718
rect 1061 704 1066 718
rect 1077 704 1082 718
rect 1140 712 1145 717
rect 1198 706 1203 725
rect 1221 706 1226 725
rect 1872 704 1877 728
rect 1895 704 1900 728
rect 1953 718 1958 721
rect 1953 704 1958 713
rect 2008 704 2013 728
rect 2031 704 2036 728
rect 2089 718 2094 721
rect 2089 704 2094 713
rect 2154 706 2159 730
rect 2177 706 2182 730
rect 2235 720 2240 723
rect 2235 706 2240 715
rect 2301 706 2306 730
rect 2324 706 2329 730
rect 2382 720 2387 723
rect 2382 706 2387 715
rect 1954 700 1958 704
rect 484 683 489 686
rect 323 660 328 678
rect 341 672 346 678
rect 1872 680 1877 699
rect 406 660 411 678
rect 323 655 411 660
rect 424 643 429 678
rect 484 669 489 678
rect 1895 680 1900 699
rect 1953 696 1958 700
rect 2090 700 2094 704
rect 2236 702 2240 706
rect 1953 686 1958 691
rect 2008 680 2013 699
rect 2031 680 2036 699
rect 2089 696 2094 700
rect 2089 686 2094 691
rect 2154 682 2159 701
rect 2177 682 2182 701
rect 2235 698 2240 702
rect 2383 702 2387 706
rect 2513 705 2518 729
rect 2536 705 2541 729
rect 2594 719 2599 722
rect 2594 705 2599 714
rect 2649 705 2654 729
rect 2672 705 2677 729
rect 2730 719 2735 722
rect 2730 705 2735 714
rect 2795 707 2800 731
rect 2818 707 2823 731
rect 2876 721 2881 724
rect 2876 707 2881 716
rect 2942 707 2947 731
rect 2965 707 2970 731
rect 3023 721 3028 724
rect 3023 707 3028 716
rect 2235 688 2240 693
rect 2301 682 2306 701
rect 2324 682 2329 701
rect 2382 698 2387 702
rect 2595 701 2599 705
rect 2382 688 2387 693
rect 2513 681 2518 700
rect 2536 681 2541 700
rect 2594 697 2599 701
rect 2731 701 2735 705
rect 2877 703 2881 707
rect 2594 687 2599 692
rect 2649 681 2654 700
rect 2672 681 2677 700
rect 2730 697 2735 701
rect 2730 687 2735 692
rect 2795 683 2800 702
rect 2818 683 2823 702
rect 2876 699 2881 703
rect 3024 703 3028 707
rect 2876 689 2881 694
rect 2942 683 2947 702
rect 2965 683 2970 702
rect 3023 699 3028 703
rect 3023 689 3028 694
rect 485 665 489 669
rect 484 661 489 665
rect 484 651 489 656
rect 1872 625 1877 639
rect 1895 625 1900 639
rect 2016 625 2021 639
rect 2039 625 2044 639
rect 2165 627 2170 641
rect 2188 627 2193 641
rect 2310 628 2315 642
rect 2333 628 2338 642
rect 1872 596 1877 620
rect 1895 596 1900 620
rect 1953 610 1958 613
rect 1953 596 1958 605
rect 2016 596 2021 620
rect 2039 596 2044 620
rect 2097 610 2102 613
rect 2097 596 2102 605
rect 2165 598 2170 622
rect 2188 598 2193 622
rect 2246 612 2251 615
rect 2246 598 2251 607
rect 2310 599 2315 623
rect 2333 599 2338 623
rect 2391 613 2396 616
rect 2391 599 2396 608
rect 1954 592 1958 596
rect 1872 572 1877 591
rect 1565 555 1570 569
rect 1588 555 1593 569
rect 1895 572 1900 591
rect 1953 588 1958 592
rect 2098 592 2102 596
rect 2247 594 2251 598
rect 2392 595 2396 599
rect 1953 578 1958 583
rect 2016 572 2021 591
rect 2039 572 2044 591
rect 2097 588 2102 592
rect 2097 578 2102 583
rect 2165 574 2170 593
rect 2188 574 2193 593
rect 2246 590 2251 594
rect 2246 580 2251 585
rect 2310 575 2315 594
rect 2333 575 2338 594
rect 2391 591 2396 595
rect 2391 581 2396 586
rect 338 521 376 522
rect 381 521 426 522
rect 338 517 426 521
rect 209 504 214 507
rect 269 504 274 507
rect 320 500 325 504
rect 338 500 343 517
rect 403 500 408 504
rect 421 500 426 517
rect 751 513 756 527
rect 774 513 779 527
rect 898 513 903 527
rect 921 513 926 527
rect 1565 526 1570 550
rect 1588 526 1593 550
rect 1644 541 1649 544
rect 1644 527 1649 536
rect 1044 511 1049 525
rect 1067 511 1072 525
rect 1180 511 1185 525
rect 1203 511 1208 525
rect 1645 523 1649 527
rect 209 490 214 499
rect 210 486 214 490
rect 209 482 214 486
rect 269 490 274 499
rect 693 498 698 501
rect 269 486 273 490
rect 269 482 274 486
rect 320 483 325 495
rect 338 491 343 495
rect 403 483 408 495
rect 421 491 426 495
rect 693 484 698 493
rect 751 484 756 508
rect 774 484 779 508
rect 840 498 845 501
rect 840 484 845 493
rect 898 484 903 508
rect 921 484 926 508
rect 986 496 991 499
rect 321 478 343 483
rect 403 478 426 483
rect 209 472 214 477
rect 269 472 274 477
rect 301 466 325 471
rect 301 458 306 466
rect 320 461 325 466
rect 338 461 343 478
rect 403 461 408 465
rect 421 461 426 478
rect 693 480 697 484
rect 693 476 698 480
rect 840 480 844 484
rect 693 466 698 471
rect 481 461 486 464
rect 751 460 756 479
rect 320 438 325 456
rect 338 450 343 456
rect 403 438 408 456
rect 320 433 408 438
rect 421 421 426 456
rect 481 447 486 456
rect 774 460 779 479
rect 840 476 845 480
rect 986 482 991 491
rect 1044 482 1049 506
rect 1067 482 1072 506
rect 1122 496 1127 499
rect 1122 482 1127 491
rect 1180 482 1185 506
rect 1203 482 1208 506
rect 1565 502 1570 521
rect 1588 502 1593 521
rect 1644 519 1649 523
rect 1644 510 1649 514
rect 840 466 845 471
rect 898 460 903 479
rect 921 460 926 479
rect 986 478 990 482
rect 986 474 991 478
rect 1122 478 1126 482
rect 986 464 991 469
rect 1044 458 1049 477
rect 1067 458 1072 477
rect 1122 474 1127 478
rect 1122 464 1127 469
rect 1180 458 1185 477
rect 1203 458 1208 477
rect 482 443 486 447
rect 481 439 486 443
rect 1564 437 1569 451
rect 1587 437 1592 451
rect 481 429 486 434
rect 742 406 747 420
rect 765 406 770 420
rect 887 405 892 419
rect 910 405 915 419
rect 684 391 689 394
rect 684 377 689 386
rect 742 377 747 401
rect 765 377 770 401
rect 1036 403 1041 417
rect 1059 403 1064 417
rect 1180 403 1185 417
rect 1203 403 1208 417
rect 1564 408 1569 432
rect 1587 408 1592 432
rect 1643 422 1648 425
rect 1643 408 1648 417
rect 829 390 834 393
rect 684 373 688 377
rect 684 369 689 373
rect 829 376 834 385
rect 887 376 892 400
rect 910 376 915 400
rect 1416 402 1421 405
rect 1454 402 1459 405
rect 1644 404 1648 408
rect 978 388 983 391
rect 829 372 833 376
rect 684 359 689 364
rect 742 353 747 372
rect 765 353 770 372
rect 829 368 834 372
rect 978 374 983 383
rect 1036 374 1041 398
rect 1059 374 1064 398
rect 1122 388 1127 391
rect 1122 374 1127 383
rect 1180 374 1185 398
rect 1203 374 1208 398
rect 1416 388 1421 397
rect 1454 388 1459 397
rect 1417 384 1421 388
rect 1455 384 1459 388
rect 1416 380 1421 384
rect 1454 380 1459 384
rect 1564 384 1569 403
rect 1587 384 1592 403
rect 1643 400 1648 404
rect 1643 390 1648 395
rect 829 358 834 363
rect 887 352 892 371
rect 910 352 915 371
rect 978 370 982 374
rect 978 366 983 370
rect 1122 370 1126 374
rect 978 356 983 361
rect 1036 350 1041 369
rect 18 331 23 334
rect 77 327 82 346
rect 93 327 98 346
rect 1059 350 1064 369
rect 1122 366 1127 370
rect 1416 370 1421 375
rect 1454 370 1459 375
rect 1122 356 1127 361
rect 1180 350 1185 369
rect 1203 350 1208 369
rect 341 336 379 337
rect 384 336 429 337
rect 341 332 429 336
rect 1563 333 1568 347
rect 1586 333 1591 347
rect 109 327 114 331
rect 125 327 130 331
rect 18 317 23 326
rect 18 313 22 317
rect 18 309 23 313
rect 18 299 23 304
rect 77 293 82 322
rect 93 293 98 322
rect 109 293 114 322
rect 125 293 130 322
rect 212 319 217 322
rect 272 319 277 322
rect 323 315 328 319
rect 341 315 346 332
rect 406 315 411 319
rect 424 315 429 332
rect 212 305 217 314
rect 213 301 217 305
rect 212 297 217 301
rect 272 305 277 314
rect 272 301 276 305
rect 272 297 277 301
rect 323 298 328 310
rect 341 306 346 310
rect 406 298 411 310
rect 424 306 429 310
rect 1563 304 1568 328
rect 1586 304 1591 328
rect 1644 318 1649 321
rect 1644 304 1649 313
rect 1645 300 1649 304
rect 324 293 346 298
rect 406 293 429 298
rect 77 281 82 288
rect 93 281 98 288
rect 109 271 114 288
rect 125 271 130 288
rect 212 287 217 292
rect 272 287 277 292
rect 304 281 328 286
rect 304 273 309 281
rect 323 276 328 281
rect 341 276 346 293
rect 406 276 411 280
rect 424 276 429 293
rect 1563 280 1568 299
rect 484 276 489 279
rect 323 253 328 271
rect 341 265 346 271
rect 1586 280 1591 299
rect 1644 296 1649 300
rect 1644 286 1649 291
rect 406 253 411 271
rect 323 248 411 253
rect 424 236 429 271
rect 484 262 489 271
rect 485 258 489 262
rect 484 254 489 258
rect 484 244 489 249
rect 1563 237 1568 251
rect 1586 237 1591 251
rect 1563 208 1568 232
rect 1586 208 1591 232
rect 1643 222 1648 225
rect 1643 208 1648 217
rect 1644 204 1648 208
rect 1563 184 1568 203
rect 1586 184 1591 203
rect 1643 200 1648 204
rect 1643 190 1648 195
rect 341 161 379 162
rect 384 161 429 162
rect 341 157 429 161
rect 212 144 217 147
rect 272 144 277 147
rect 323 140 328 144
rect 341 140 346 157
rect 406 140 411 144
rect 424 140 429 157
rect 212 130 217 139
rect 213 126 217 130
rect 212 122 217 126
rect 272 130 277 139
rect 272 126 276 130
rect 272 122 277 126
rect 323 123 328 135
rect 341 131 346 135
rect 406 123 411 135
rect 424 131 429 135
rect 324 118 346 123
rect 406 118 429 123
rect 212 112 217 117
rect 272 112 277 117
rect 304 106 328 111
rect 304 98 309 106
rect 323 101 328 106
rect 341 101 346 118
rect 406 101 411 105
rect 424 101 429 118
rect 484 101 489 104
rect 323 78 328 96
rect 341 90 346 96
rect 406 78 411 96
rect 323 73 411 78
rect 424 61 429 96
rect 484 87 489 96
rect 485 83 489 87
rect 484 79 489 83
rect 484 69 489 74
<< polycontact >>
rect 882 1029 887 1033
rect 936 1003 941 1009
rect 959 1003 964 1009
rect 774 947 779 951
rect 831 948 836 952
rect 669 902 674 909
rect 685 902 690 909
rect 701 902 706 909
rect 717 903 722 910
rect 722 777 727 782
rect 738 777 744 783
rect 883 777 889 784
rect 899 777 905 784
rect 931 777 937 783
rect 1060 779 1067 785
rect 379 743 384 748
rect 639 744 644 748
rect 1075 777 1085 785
rect 828 744 833 748
rect 986 744 991 748
rect 208 708 213 712
rect 1144 726 1149 730
rect 276 708 281 712
rect 319 700 324 705
rect 915 696 922 702
rect 1043 696 1051 703
rect 1198 700 1203 706
rect 1221 700 1226 706
rect 1949 700 1954 704
rect 304 675 309 680
rect 1872 674 1877 680
rect 2085 700 2090 704
rect 2231 702 2236 706
rect 1895 674 1900 680
rect 2008 674 2013 680
rect 2031 674 2036 680
rect 2154 676 2159 682
rect 2378 702 2383 706
rect 2177 676 2182 682
rect 2301 676 2306 682
rect 2590 701 2595 705
rect 2324 676 2329 682
rect 2513 675 2518 681
rect 2726 701 2731 705
rect 2872 703 2877 707
rect 2536 675 2541 681
rect 2649 675 2654 681
rect 2672 675 2677 681
rect 2795 677 2800 683
rect 3019 703 3024 707
rect 2818 677 2823 683
rect 2942 677 2947 683
rect 2965 677 2970 683
rect 480 665 485 669
rect 424 638 429 643
rect 1949 592 1954 596
rect 1872 566 1877 572
rect 2093 592 2098 596
rect 2242 594 2247 598
rect 2387 595 2392 599
rect 1895 566 1900 572
rect 2016 566 2021 572
rect 2039 566 2044 572
rect 2165 568 2170 574
rect 2188 568 2193 574
rect 2310 569 2315 575
rect 2333 569 2338 575
rect 376 521 381 526
rect 1640 523 1645 527
rect 205 486 210 490
rect 273 486 278 490
rect 316 478 321 483
rect 301 453 306 458
rect 697 480 702 484
rect 844 480 849 484
rect 751 454 756 460
rect 1565 496 1570 502
rect 1588 496 1593 502
rect 774 454 779 460
rect 898 454 903 460
rect 990 478 995 482
rect 1126 478 1131 482
rect 921 454 926 460
rect 1044 452 1049 458
rect 1067 452 1072 458
rect 1180 452 1185 458
rect 1203 452 1208 458
rect 477 443 482 447
rect 421 416 426 421
rect 688 373 693 377
rect 1639 404 1644 408
rect 833 372 838 376
rect 77 346 83 353
rect 93 346 99 353
rect 742 347 747 353
rect 1412 384 1417 388
rect 1450 384 1455 388
rect 1564 378 1569 384
rect 1587 378 1592 384
rect 765 347 770 353
rect 887 346 892 352
rect 982 370 987 374
rect 1126 370 1131 374
rect 910 346 915 352
rect 1036 344 1041 350
rect 1059 344 1064 350
rect 1180 344 1185 350
rect 1203 344 1208 350
rect 379 336 384 341
rect 22 313 27 317
rect 208 301 213 305
rect 276 301 281 305
rect 1640 300 1645 304
rect 319 293 324 298
rect 109 265 116 271
rect 125 265 132 271
rect 304 268 309 273
rect 1563 274 1568 280
rect 1586 274 1591 280
rect 480 258 485 262
rect 424 231 429 236
rect 1639 204 1644 208
rect 1563 178 1568 184
rect 1586 178 1591 184
rect 379 161 384 166
rect 208 126 213 130
rect 276 126 281 130
rect 319 118 324 123
rect 304 93 309 98
rect 480 83 485 87
rect 424 56 429 61
<< metal1 >>
rect 904 1073 932 1074
rect 904 1070 990 1073
rect 904 1060 908 1070
rect 929 1069 990 1070
rect 929 1068 980 1069
rect 929 1062 934 1068
rect 966 1062 971 1068
rect 904 1059 909 1060
rect 861 1054 909 1059
rect 975 1062 980 1068
rect 885 1047 890 1054
rect 897 1047 902 1054
rect 947 1047 952 1057
rect 947 1043 957 1047
rect 870 1033 875 1042
rect 953 1039 957 1043
rect 916 1036 957 1039
rect 916 1033 919 1036
rect 953 1033 957 1036
rect 859 1029 875 1033
rect 887 1029 919 1033
rect 870 1025 875 1029
rect 927 1028 929 1031
rect 885 1016 890 1020
rect 927 1017 930 1028
rect 944 1025 947 1028
rect 971 1017 974 1031
rect 859 1011 895 1016
rect 859 1010 866 1011
rect 927 1012 974 1017
rect 859 989 864 1010
rect 936 1002 941 1003
rect 959 987 964 1003
rect 950 984 964 987
rect 809 977 857 978
rect 985 977 990 1069
rect 1247 977 1270 978
rect 647 974 1271 977
rect 647 973 1262 974
rect 647 972 800 973
rect 661 961 666 972
rect 737 961 742 972
rect 759 965 764 972
rect 771 965 776 972
rect 816 966 821 973
rect 828 966 833 973
rect 725 934 730 956
rect 786 951 791 960
rect 843 952 848 961
rect 944 952 948 960
rect 795 951 831 952
rect 756 947 774 951
rect 786 948 831 951
rect 843 948 948 952
rect 786 947 829 948
rect 756 934 759 947
rect 786 943 791 947
rect 843 944 848 948
rect 771 934 776 938
rect 828 935 833 939
rect 819 934 858 935
rect 677 930 759 934
rect 762 930 882 934
rect 677 925 682 930
rect 709 925 714 930
rect 762 929 801 930
rect 889 930 1181 934
rect 661 916 666 920
rect 693 917 698 920
rect 725 917 730 920
rect 762 917 767 929
rect 693 916 767 917
rect 661 913 767 916
rect 669 900 674 902
rect 685 898 690 902
rect 685 885 689 898
rect 701 897 706 902
rect 722 903 866 904
rect 717 899 866 903
rect 1178 903 1181 930
rect 1266 921 1271 974
rect 685 882 795 885
rect 292 873 934 875
rect 292 872 935 873
rect 292 808 295 872
rect 655 849 660 864
rect 796 849 800 864
rect 931 851 935 872
rect 141 805 295 808
rect 178 804 295 805
rect 578 837 585 840
rect 928 837 952 838
rect 578 834 1066 837
rect 94 782 186 784
rect 93 777 186 782
rect 76 354 82 763
rect 77 353 82 354
rect 93 544 99 777
rect 460 763 461 769
rect 475 763 554 769
rect 379 750 530 755
rect 178 746 372 750
rect 178 712 183 746
rect 193 734 356 738
rect 193 733 308 734
rect 193 726 198 733
rect 205 726 210 733
rect 279 726 284 733
rect 220 712 225 721
rect 291 726 296 733
rect 303 722 308 733
rect 178 709 208 712
rect 204 708 208 709
rect 220 708 229 712
rect 264 712 269 721
rect 315 722 320 734
rect 238 708 269 712
rect 281 708 287 712
rect 220 704 225 708
rect 205 695 210 699
rect 196 690 227 695
rect 238 644 242 708
rect 264 704 269 708
rect 294 708 302 712
rect 298 705 302 708
rect 349 711 354 717
rect 367 711 372 746
rect 379 748 384 750
rect 398 728 451 734
rect 398 722 403 728
rect 432 711 437 717
rect 349 706 437 711
rect 298 700 319 705
rect 279 695 284 699
rect 255 690 293 695
rect 283 653 288 690
rect 349 683 354 706
rect 304 672 309 675
rect 383 682 389 695
rect 315 653 320 678
rect 398 683 403 693
rect 432 683 437 706
rect 446 653 451 728
rect 463 690 506 695
rect 465 683 470 690
rect 477 683 482 690
rect 492 670 497 678
rect 511 670 516 750
rect 548 680 554 763
rect 578 715 585 834
rect 717 824 736 829
rect 607 698 611 823
rect 655 786 660 823
rect 717 788 725 824
rect 796 788 800 826
rect 853 794 889 801
rect 717 787 743 788
rect 717 785 744 787
rect 736 783 744 785
rect 690 777 722 782
rect 736 781 738 783
rect 882 785 888 794
rect 883 784 888 785
rect 899 784 904 789
rect 931 783 935 825
rect 1061 785 1066 834
rect 1077 803 1081 853
rect 1178 795 1182 903
rect 1265 901 1271 921
rect 1077 785 1081 792
rect 617 770 1130 774
rect 1265 772 1270 901
rect 1248 771 1349 772
rect 618 769 666 770
rect 642 762 647 769
rect 654 762 659 769
rect 698 758 703 770
rect 730 758 735 770
rect 762 758 767 770
rect 807 769 855 770
rect 627 748 632 757
rect 831 762 836 769
rect 682 750 687 753
rect 714 750 719 753
rect 682 749 719 750
rect 746 749 751 753
rect 622 744 632 748
rect 644 745 668 748
rect 644 744 659 745
rect 627 740 632 744
rect 642 731 647 735
rect 664 736 668 745
rect 682 745 751 749
rect 796 748 800 758
rect 843 762 848 769
rect 863 758 868 770
rect 816 748 821 757
rect 875 758 880 770
rect 907 758 912 770
rect 939 758 944 770
rect 965 769 1130 770
rect 989 762 994 769
rect 1001 762 1006 769
rect 1027 757 1032 769
rect 1053 757 1058 769
rect 1085 757 1090 769
rect 891 750 896 753
rect 876 749 896 750
rect 923 749 928 753
rect 682 736 687 745
rect 796 744 821 748
rect 833 744 852 748
rect 664 731 687 736
rect 816 740 821 744
rect 831 731 836 735
rect 848 736 852 744
rect 876 745 928 749
rect 876 736 881 745
rect 974 748 979 757
rect 1036 752 1037 757
rect 1124 756 1130 769
rect 1163 770 1194 771
rect 1241 770 1349 771
rect 1163 767 1349 770
rect 1167 756 1171 767
rect 1036 749 1042 752
rect 1069 749 1074 752
rect 1123 751 1171 756
rect 1191 765 1242 767
rect 1248 766 1349 767
rect 1191 759 1196 765
rect 1228 759 1233 765
rect 1237 759 1242 765
rect 967 744 979 748
rect 991 744 1017 748
rect 1036 744 1074 749
rect 1147 744 1152 751
rect 848 731 881 736
rect 974 740 979 744
rect 989 731 994 735
rect 1013 731 1017 744
rect 1034 731 1039 744
rect 1159 744 1164 751
rect 1209 744 1214 754
rect 1209 740 1219 744
rect 617 726 656 731
rect 651 710 656 726
rect 682 724 687 731
rect 806 726 845 731
rect 762 712 767 719
rect 840 712 845 726
rect 876 724 881 731
rect 963 726 1009 731
rect 1013 726 1039 731
rect 762 710 845 712
rect 939 717 944 719
rect 964 717 970 726
rect 939 714 970 717
rect 1005 725 1009 726
rect 939 713 949 714
rect 939 710 944 713
rect 651 707 944 710
rect 1005 711 1010 725
rect 1034 723 1039 726
rect 1132 730 1137 739
rect 1215 736 1219 740
rect 1178 733 1219 736
rect 1178 730 1181 733
rect 1215 730 1219 733
rect 1126 726 1137 730
rect 1149 726 1181 730
rect 1085 711 1090 718
rect 1132 722 1137 726
rect 1189 725 1191 728
rect 1147 713 1152 717
rect 1189 714 1192 725
rect 1206 722 1209 725
rect 1233 714 1236 728
rect 1121 711 1157 713
rect 1005 708 1157 711
rect 1005 707 1130 708
rect 1189 709 1236 714
rect 651 706 767 707
rect 840 706 944 707
rect 607 696 690 698
rect 607 694 695 696
rect 706 689 711 696
rect 754 693 759 696
rect 706 685 737 689
rect 548 678 683 680
rect 548 675 684 678
rect 477 665 480 669
rect 492 665 516 670
rect 492 661 497 665
rect 678 661 684 675
rect 728 674 736 685
rect 730 666 736 674
rect 753 680 762 693
rect 915 692 920 696
rect 1045 693 1049 696
rect 753 673 755 680
rect 728 665 736 666
rect 283 652 451 653
rect 477 652 482 656
rect 283 648 530 652
rect 446 647 530 648
rect 238 639 407 644
rect 402 634 407 639
rect 424 634 429 638
rect 402 629 429 634
rect 93 541 224 544
rect 93 540 99 541
rect 93 353 98 540
rect 507 533 514 599
rect 376 528 514 533
rect 175 524 369 528
rect 175 490 180 524
rect 190 512 353 516
rect 190 511 305 512
rect 190 504 195 511
rect 202 504 207 511
rect 276 504 281 511
rect 217 490 222 499
rect 288 504 293 511
rect 300 500 305 511
rect 175 487 205 490
rect 201 486 205 487
rect 217 486 226 490
rect 261 490 266 499
rect 312 500 317 512
rect 235 486 266 490
rect 278 488 299 490
rect 278 486 286 488
rect 217 482 222 486
rect 202 473 207 477
rect 193 468 224 473
rect 235 422 239 486
rect 261 482 266 486
rect 292 486 299 488
rect 295 483 299 486
rect 346 489 351 495
rect 364 489 369 524
rect 376 526 381 528
rect 395 506 448 512
rect 395 500 400 506
rect 429 489 434 495
rect 346 484 434 489
rect 295 478 316 483
rect 276 473 281 477
rect 252 468 290 473
rect 280 431 285 468
rect 346 461 351 484
rect 395 478 398 481
rect 388 473 403 478
rect 301 450 306 453
rect 380 462 385 473
rect 395 461 400 473
rect 429 461 434 484
rect 312 431 317 456
rect 443 431 448 506
rect 460 468 503 473
rect 462 461 467 468
rect 474 461 479 468
rect 489 448 494 456
rect 508 448 513 528
rect 474 443 477 447
rect 489 443 513 448
rect 523 465 529 647
rect 548 610 557 648
rect 677 655 684 661
rect 570 596 577 647
rect 620 623 621 630
rect 620 566 627 623
rect 552 558 628 566
rect 677 558 683 655
rect 739 617 748 642
rect 914 638 920 692
rect 1044 630 1049 693
rect 1121 685 1130 707
rect 1198 699 1203 700
rect 1221 699 1226 700
rect 1122 676 1130 685
rect 1122 675 1322 676
rect 1122 673 1325 675
rect 1318 665 1325 673
rect 739 611 1109 617
rect 789 579 815 585
rect 1102 577 1109 611
rect 727 562 958 566
rect 1319 561 1323 665
rect 676 553 683 558
rect 585 532 651 539
rect 677 510 683 553
rect 716 524 747 525
rect 794 524 894 525
rect 716 523 942 524
rect 716 522 1040 523
rect 1145 522 1176 523
rect 1343 522 1347 766
rect 1676 767 1991 771
rect 1855 766 1991 767
rect 2071 764 2076 807
rect 2118 797 2618 802
rect 2118 777 2124 797
rect 2071 760 2132 764
rect 2188 763 2193 778
rect 2271 774 2766 780
rect 2188 760 2281 763
rect 1693 744 1700 749
rect 2827 747 2927 748
rect 2974 747 3005 748
rect 2186 746 2286 747
rect 2333 746 2364 747
rect 2779 746 3005 747
rect 2132 745 2364 746
rect 2545 745 2576 746
rect 2681 745 3005 746
rect 1904 744 1935 745
rect 2040 744 2364 745
rect 2490 744 3005 745
rect 1693 743 2830 744
rect 1693 741 2189 743
rect 1693 739 1907 741
rect 1471 566 1476 568
rect 1693 567 1700 739
rect 1835 738 1862 739
rect 1835 638 1843 738
rect 1856 733 1861 738
rect 1865 733 1870 739
rect 1902 733 1907 739
rect 1927 740 2043 741
rect 1927 730 1931 740
rect 1992 739 2043 740
rect 1992 733 1997 739
rect 1884 718 1889 728
rect 1927 725 1975 730
rect 2001 733 2006 739
rect 2038 733 2043 739
rect 2063 730 2067 741
rect 2139 735 2143 741
rect 2147 735 2152 741
rect 2184 735 2189 741
rect 2209 732 2213 743
rect 2285 741 2336 743
rect 2285 735 2290 741
rect 1879 714 1889 718
rect 1934 718 1939 725
rect 1879 710 1883 714
rect 1946 718 1951 725
rect 2020 718 2025 728
rect 2063 725 2111 730
rect 1879 707 1920 710
rect 1879 704 1883 707
rect 1917 704 1920 707
rect 1961 704 1966 713
rect 2015 714 2025 718
rect 2070 718 2075 725
rect 2015 710 2019 714
rect 2082 718 2087 725
rect 2166 720 2171 730
rect 2209 727 2257 732
rect 2294 735 2299 741
rect 2331 735 2336 741
rect 2356 742 2830 743
rect 2356 740 2548 742
rect 2356 732 2360 740
rect 2490 739 2503 740
rect 2497 734 2502 739
rect 2015 707 2056 710
rect 1862 688 1865 702
rect 1907 699 1909 702
rect 1917 700 1949 704
rect 1961 700 1980 704
rect 1889 696 1892 699
rect 1906 688 1909 699
rect 1961 696 1966 700
rect 2015 704 2019 707
rect 2053 704 2056 707
rect 2097 704 2102 713
rect 2161 716 2171 720
rect 2216 720 2221 727
rect 2161 712 2165 716
rect 2228 720 2233 727
rect 2313 720 2318 730
rect 2356 727 2404 732
rect 2506 734 2511 740
rect 2543 734 2548 740
rect 2568 741 2684 742
rect 2568 731 2572 741
rect 2633 740 2684 741
rect 2633 734 2638 740
rect 2161 709 2202 712
rect 2161 706 2165 709
rect 2199 706 2202 709
rect 2243 706 2248 715
rect 2308 716 2318 720
rect 2363 720 2368 727
rect 2308 712 2312 716
rect 2375 720 2380 727
rect 2525 719 2530 729
rect 2568 726 2616 731
rect 2642 734 2647 740
rect 2679 734 2684 740
rect 2704 731 2708 742
rect 2779 736 2784 742
rect 2788 736 2793 742
rect 2825 736 2830 742
rect 2850 733 2854 744
rect 2926 742 2977 744
rect 2926 736 2931 742
rect 2308 709 2349 712
rect 1862 683 1909 688
rect 1946 687 1951 691
rect 1998 688 2001 702
rect 2043 699 2045 702
rect 2053 700 2085 704
rect 2097 700 2118 704
rect 2025 696 2028 699
rect 2042 688 2045 699
rect 2097 696 2102 700
rect 1941 682 1976 687
rect 1998 683 2045 688
rect 1872 673 1877 674
rect 1895 673 1900 674
rect 1972 661 1976 682
rect 2082 687 2087 691
rect 2144 690 2147 704
rect 2189 701 2191 704
rect 2199 702 2231 706
rect 2243 702 2264 706
rect 2171 698 2174 701
rect 2188 690 2191 701
rect 2243 698 2248 702
rect 2308 706 2312 709
rect 2346 706 2349 709
rect 2390 706 2395 715
rect 2520 715 2530 719
rect 2575 719 2580 726
rect 2520 711 2524 715
rect 2587 719 2592 726
rect 2661 719 2666 729
rect 2704 726 2752 731
rect 2520 708 2561 711
rect 2077 686 2112 687
rect 2077 682 2125 686
rect 2144 685 2191 690
rect 2228 689 2233 693
rect 2291 690 2294 704
rect 2336 701 2338 704
rect 2346 702 2378 706
rect 2390 702 2420 706
rect 2318 698 2321 701
rect 2335 690 2338 701
rect 2390 698 2395 702
rect 2520 705 2524 708
rect 2558 705 2561 708
rect 2602 705 2607 714
rect 2656 715 2666 719
rect 2711 719 2716 726
rect 2656 711 2660 715
rect 2723 719 2728 726
rect 2807 721 2812 731
rect 2850 728 2898 733
rect 2935 736 2940 742
rect 2972 736 2977 742
rect 2997 733 3001 744
rect 2656 708 2697 711
rect 2656 705 2660 708
rect 2694 705 2697 708
rect 2738 705 2743 714
rect 2802 717 2812 721
rect 2857 721 2862 728
rect 2802 713 2806 717
rect 2869 721 2874 728
rect 2954 721 2959 731
rect 2997 728 3045 733
rect 2802 710 2843 713
rect 2802 707 2806 710
rect 2840 707 2843 710
rect 2884 707 2889 716
rect 2949 717 2959 721
rect 3004 721 3009 728
rect 2949 713 2953 717
rect 3016 721 3021 728
rect 2949 710 2990 713
rect 2949 707 2953 710
rect 2987 707 2990 710
rect 3031 707 3036 716
rect 2223 684 2261 689
rect 2291 685 2338 690
rect 2106 681 2125 682
rect 2008 673 2013 674
rect 2031 673 2036 674
rect 2116 661 2123 681
rect 2154 675 2159 676
rect 2177 675 2182 676
rect 2252 661 2261 684
rect 2375 689 2380 693
rect 2503 689 2506 703
rect 2548 700 2550 703
rect 2558 701 2590 705
rect 2602 701 2610 705
rect 2530 697 2533 700
rect 2547 689 2550 700
rect 2602 697 2607 701
rect 2370 684 2406 689
rect 2503 684 2550 689
rect 2301 675 2306 676
rect 2324 675 2329 676
rect 2397 661 2406 684
rect 2587 688 2592 692
rect 2639 689 2642 703
rect 2684 700 2686 703
rect 2694 701 2726 705
rect 2738 701 2746 705
rect 2666 697 2669 700
rect 2683 689 2686 700
rect 2738 697 2743 701
rect 2582 683 2617 688
rect 2639 684 2686 689
rect 2513 674 2518 675
rect 2536 674 2541 675
rect 2613 662 2617 683
rect 2723 688 2728 692
rect 2785 691 2788 705
rect 2830 702 2832 705
rect 2840 703 2872 707
rect 2884 703 2892 707
rect 2812 699 2815 702
rect 2829 691 2832 702
rect 2884 699 2889 703
rect 2718 687 2753 688
rect 2718 683 2766 687
rect 2785 686 2832 691
rect 2869 690 2874 694
rect 2932 691 2935 705
rect 2977 702 2979 705
rect 2987 703 3019 707
rect 3031 703 3039 707
rect 2959 699 2962 702
rect 2976 691 2979 702
rect 3031 699 3036 703
rect 2864 685 2902 690
rect 2932 686 2979 691
rect 2747 682 2766 683
rect 2649 674 2654 675
rect 2672 674 2677 675
rect 2757 662 2764 682
rect 2795 676 2800 677
rect 2818 676 2823 677
rect 2893 662 2902 685
rect 3016 690 3021 694
rect 3011 685 3047 690
rect 2942 676 2947 677
rect 2965 676 2970 677
rect 3038 662 3047 685
rect 2425 661 2433 662
rect 1972 655 2433 661
rect 2613 657 3048 662
rect 2613 656 3023 657
rect 2425 644 2433 655
rect 2634 644 2643 656
rect 2342 639 2373 640
rect 2197 638 2373 639
rect 1835 636 1865 638
rect 2073 637 2373 638
rect 1904 636 1935 637
rect 2048 636 2373 637
rect 2424 636 2643 644
rect 1835 635 2345 636
rect 1835 633 2200 635
rect 2209 634 2345 635
rect 1835 631 1907 633
rect 1926 631 2051 633
rect 1856 625 1861 631
rect 1865 625 1870 631
rect 1902 625 1907 631
rect 1927 622 1931 631
rect 2000 625 2005 631
rect 1884 610 1889 620
rect 1927 617 1975 622
rect 2009 625 2014 631
rect 2046 625 2051 631
rect 2071 622 2075 633
rect 2149 627 2154 633
rect 2158 627 2163 633
rect 2195 627 2200 633
rect 2220 624 2224 634
rect 2294 628 2299 634
rect 1879 606 1889 610
rect 1934 610 1939 617
rect 1879 602 1883 606
rect 1946 610 1951 617
rect 2028 610 2033 620
rect 2071 617 2119 622
rect 1879 599 1920 602
rect 1879 596 1883 599
rect 1917 596 1920 599
rect 1961 596 1966 605
rect 2023 606 2033 610
rect 2078 610 2083 617
rect 2023 602 2027 606
rect 2090 610 2095 617
rect 2177 612 2182 622
rect 2220 619 2268 624
rect 2303 628 2308 634
rect 2340 628 2345 634
rect 2365 625 2369 636
rect 2023 599 2064 602
rect 1862 580 1865 594
rect 1907 591 1909 594
rect 1917 592 1949 596
rect 1961 592 1993 596
rect 1889 588 1892 591
rect 1906 580 1909 591
rect 1961 588 1966 592
rect 2023 596 2027 599
rect 2061 596 2064 599
rect 2105 596 2110 605
rect 2172 608 2182 612
rect 2227 612 2232 619
rect 2172 604 2176 608
rect 2239 612 2244 619
rect 2322 613 2327 623
rect 2365 620 2413 625
rect 2172 601 2213 604
rect 2172 598 2176 601
rect 2210 598 2213 601
rect 2254 598 2259 607
rect 2317 609 2327 613
rect 2372 613 2377 620
rect 2317 605 2321 609
rect 2384 613 2389 620
rect 2317 602 2358 605
rect 2317 599 2321 602
rect 2355 599 2358 602
rect 2399 599 2404 608
rect 1862 575 1909 580
rect 1946 579 1951 583
rect 2006 580 2009 594
rect 2051 591 2053 594
rect 2061 592 2093 596
rect 2105 592 2133 596
rect 2033 588 2036 591
rect 2050 580 2053 591
rect 2105 588 2110 592
rect 1941 574 1976 579
rect 2006 575 2053 580
rect 1597 566 1700 567
rect 1471 563 1701 566
rect 1471 562 1600 563
rect 1471 522 1476 562
rect 1549 561 1600 562
rect 1549 555 1554 561
rect 1558 555 1563 561
rect 1595 555 1600 561
rect 1620 553 1624 563
rect 1693 553 1701 563
rect 1872 565 1877 566
rect 1895 565 1900 566
rect 1577 540 1582 550
rect 1618 548 1701 553
rect 1572 536 1582 540
rect 1625 541 1630 548
rect 1637 541 1642 548
rect 1572 532 1576 536
rect 1572 529 1613 532
rect 1572 526 1576 529
rect 1610 526 1613 529
rect 1652 527 1657 536
rect 1693 528 1701 548
rect 1617 526 1640 527
rect 716 521 1476 522
rect 720 510 724 521
rect 676 505 724 510
rect 744 519 795 521
rect 744 513 749 519
rect 781 513 786 519
rect 790 513 795 519
rect 867 510 871 521
rect 700 498 705 505
rect 712 498 717 505
rect 762 498 767 508
rect 823 505 871 510
rect 891 519 1476 521
rect 891 513 896 519
rect 928 513 933 519
rect 937 513 942 519
rect 1013 508 1017 519
rect 847 498 852 505
rect 762 494 772 498
rect 685 484 690 493
rect 768 490 772 494
rect 731 487 772 490
rect 731 484 734 487
rect 768 484 772 487
rect 859 498 864 505
rect 909 498 914 508
rect 969 503 1017 508
rect 1037 518 1153 519
rect 1037 517 1088 518
rect 1037 511 1042 517
rect 1074 511 1079 517
rect 1083 511 1088 517
rect 1149 508 1153 518
rect 909 494 919 498
rect 993 496 998 503
rect 667 480 690 484
rect 702 480 734 484
rect 685 476 690 480
rect 742 479 744 482
rect 700 467 705 471
rect 742 468 745 479
rect 759 476 762 479
rect 786 468 789 482
rect 832 484 837 493
rect 915 490 919 494
rect 878 487 919 490
rect 878 484 881 487
rect 915 484 919 487
rect 1005 496 1010 503
rect 1055 496 1060 506
rect 1105 503 1153 508
rect 1173 517 1476 519
rect 1173 511 1178 517
rect 1210 511 1215 517
rect 1218 516 1476 517
rect 1219 511 1224 516
rect 1129 496 1134 503
rect 1055 492 1065 496
rect 821 481 837 484
rect 819 480 837 481
rect 849 480 881 484
rect 832 476 837 480
rect 889 479 891 482
rect 674 465 710 467
rect 523 462 710 465
rect 523 460 683 462
rect 742 463 789 468
rect 847 467 852 471
rect 889 468 892 479
rect 906 476 909 479
rect 933 468 936 482
rect 978 482 983 491
rect 1061 488 1065 492
rect 1024 485 1065 488
rect 1024 482 1027 485
rect 1061 482 1065 485
rect 1141 496 1146 503
rect 1191 496 1196 506
rect 1191 492 1201 496
rect 1114 482 1119 491
rect 1197 488 1201 492
rect 1160 485 1201 488
rect 1160 482 1163 485
rect 1197 482 1201 485
rect 966 478 983 482
rect 995 478 1027 482
rect 978 474 983 478
rect 1035 477 1037 480
rect 1104 481 1119 482
rect 819 462 857 467
rect 489 439 494 443
rect 280 430 448 431
rect 474 430 479 434
rect 523 430 529 460
rect 280 426 529 430
rect 443 425 529 426
rect 235 417 404 422
rect 399 412 404 417
rect 421 412 426 416
rect 160 401 198 405
rect 399 407 426 412
rect 160 400 202 401
rect 483 348 488 360
rect 144 343 149 348
rect 379 343 516 348
rect 1 339 149 343
rect 153 339 372 343
rect 1 338 49 339
rect 25 331 30 338
rect 37 331 42 338
rect 57 327 62 339
rect 10 317 15 326
rect 69 327 74 339
rect 101 327 106 339
rect 133 327 138 339
rect 85 319 90 322
rect 70 318 90 319
rect 117 318 122 322
rect 3 313 15 317
rect 27 313 46 317
rect 10 309 15 313
rect 25 300 30 304
rect 42 305 46 313
rect 70 314 122 318
rect 70 305 75 314
rect 42 300 45 305
rect 50 300 75 305
rect 153 305 158 339
rect 168 327 356 331
rect 168 326 308 327
rect 168 319 173 326
rect 205 319 210 326
rect 279 319 284 326
rect 220 305 225 314
rect 291 319 296 326
rect 303 315 308 326
rect 264 305 269 314
rect 315 315 320 327
rect 153 302 208 305
rect 204 301 208 302
rect 220 301 228 305
rect 0 295 39 300
rect 34 279 39 295
rect 70 293 75 300
rect 220 297 225 301
rect 238 301 269 305
rect 281 303 302 305
rect 281 301 288 303
rect 205 288 210 292
rect 133 286 138 288
rect 171 286 227 288
rect 133 283 227 286
rect 133 282 175 283
rect 133 279 138 282
rect 34 275 138 279
rect 153 268 186 271
rect 109 249 114 265
rect 125 260 130 265
rect 125 256 226 260
rect 109 245 143 249
rect 238 237 242 301
rect 264 297 269 301
rect 293 301 302 303
rect 298 298 302 301
rect 349 304 354 310
rect 367 304 372 339
rect 379 341 384 343
rect 398 321 451 327
rect 398 315 403 321
rect 432 304 437 310
rect 349 299 437 304
rect 298 293 319 298
rect 279 288 284 292
rect 255 283 293 288
rect 283 246 288 283
rect 349 276 354 299
rect 398 293 401 296
rect 304 265 309 268
rect 391 288 406 293
rect 383 275 388 288
rect 315 246 320 271
rect 398 276 403 288
rect 432 276 437 299
rect 446 246 451 321
rect 463 283 506 288
rect 465 276 470 283
rect 477 276 482 283
rect 492 263 497 271
rect 511 263 516 343
rect 477 258 480 262
rect 492 258 516 263
rect 492 254 497 258
rect 283 245 451 246
rect 477 245 482 249
rect 523 245 529 425
rect 541 432 542 441
rect 647 439 655 440
rect 674 439 683 460
rect 751 453 756 454
rect 774 453 779 454
rect 819 439 828 462
rect 889 463 936 468
rect 993 465 998 469
rect 1035 466 1038 477
rect 1052 474 1055 477
rect 1079 466 1082 480
rect 1109 478 1119 481
rect 1131 478 1163 482
rect 1114 474 1119 478
rect 1171 477 1173 480
rect 968 464 1003 465
rect 955 460 1003 464
rect 898 453 903 454
rect 955 459 974 460
rect 1035 461 1082 466
rect 1129 465 1134 469
rect 1171 466 1174 477
rect 1188 474 1191 477
rect 1215 466 1218 480
rect 1104 460 1139 465
rect 921 453 926 454
rect 957 439 964 459
rect 1044 451 1049 452
rect 1067 451 1072 452
rect 1104 439 1108 460
rect 1171 461 1218 466
rect 1180 451 1185 452
rect 1203 451 1208 452
rect 541 389 548 432
rect 575 355 581 438
rect 647 433 1108 439
rect 545 349 581 355
rect 618 324 620 333
rect 618 256 627 324
rect 283 241 531 245
rect 446 240 531 241
rect 238 232 407 237
rect 402 227 407 232
rect 424 227 429 231
rect 402 222 429 227
rect 502 203 506 225
rect 379 168 510 173
rect 178 164 372 168
rect 178 130 183 164
rect 193 152 356 156
rect 193 151 308 152
rect 193 144 198 151
rect 205 144 210 151
rect 279 144 284 151
rect 220 130 225 139
rect 291 144 296 151
rect 303 140 308 151
rect 264 130 269 139
rect 315 140 320 152
rect 178 127 208 130
rect 204 126 208 127
rect 220 126 228 130
rect 220 122 225 126
rect 238 126 269 130
rect 281 128 302 130
rect 281 126 288 128
rect 205 113 210 117
rect 196 108 227 113
rect 238 62 242 126
rect 264 122 269 126
rect 294 126 302 128
rect 298 123 302 126
rect 349 129 354 135
rect 367 129 372 164
rect 379 166 384 168
rect 398 146 451 152
rect 398 140 403 146
rect 432 129 437 135
rect 349 124 437 129
rect 298 118 319 123
rect 279 113 284 117
rect 255 108 293 113
rect 283 71 288 108
rect 349 101 354 124
rect 398 118 401 121
rect 388 113 406 118
rect 304 90 309 93
rect 379 101 386 113
rect 398 101 403 113
rect 379 96 383 101
rect 432 101 437 124
rect 315 71 320 96
rect 446 71 451 146
rect 463 108 506 113
rect 465 101 470 108
rect 477 101 482 108
rect 492 88 497 96
rect 511 88 516 168
rect 477 83 480 87
rect 492 83 516 88
rect 492 79 497 83
rect 283 70 451 71
rect 477 70 482 74
rect 523 70 529 240
rect 617 172 627 256
rect 617 107 626 172
rect 283 66 529 70
rect 446 65 529 66
rect 238 57 407 62
rect 402 52 407 57
rect 424 52 429 56
rect 402 47 429 52
rect 476 29 483 38
rect 635 29 641 373
rect 647 327 655 433
rect 707 417 738 418
rect 707 416 883 417
rect 1237 416 1245 516
rect 707 415 1007 416
rect 707 414 1032 415
rect 1145 414 1176 415
rect 1215 414 1245 416
rect 1471 414 1476 516
rect 1555 510 1558 524
rect 1600 521 1602 524
rect 1610 523 1640 526
rect 1652 523 1660 527
rect 1610 522 1637 523
rect 1582 518 1585 521
rect 1599 510 1602 521
rect 1652 519 1657 523
rect 1694 523 1700 528
rect 1834 523 1837 553
rect 1968 550 1977 574
rect 2090 579 2095 583
rect 2155 582 2158 596
rect 2200 593 2202 596
rect 2210 594 2242 598
rect 2254 594 2282 598
rect 2182 590 2185 593
rect 2199 582 2202 593
rect 2254 590 2259 594
rect 2085 574 2126 579
rect 2155 577 2202 582
rect 2239 581 2244 585
rect 2300 583 2303 597
rect 2345 594 2347 597
rect 2355 595 2387 599
rect 2399 595 2407 599
rect 2327 591 2330 594
rect 2344 583 2347 594
rect 2399 591 2404 595
rect 2234 576 2269 581
rect 2300 578 2347 583
rect 2384 582 2389 586
rect 2408 582 2415 583
rect 2379 577 2415 582
rect 2016 565 2021 566
rect 2039 565 2044 566
rect 2118 550 2125 574
rect 2165 567 2170 568
rect 2188 567 2193 568
rect 2262 550 2269 576
rect 2310 567 2315 569
rect 2333 568 2338 569
rect 2408 550 2415 577
rect 1968 549 2415 550
rect 2425 549 2433 636
rect 2634 635 2643 636
rect 1968 544 2433 549
rect 1637 510 1642 514
rect 1555 505 1602 510
rect 1634 505 1656 510
rect 1649 504 1656 505
rect 711 403 715 414
rect 667 398 715 403
rect 735 413 1245 414
rect 735 412 871 413
rect 735 406 740 412
rect 772 406 777 412
rect 781 406 786 412
rect 856 402 860 412
rect 691 391 696 398
rect 703 391 708 398
rect 753 391 758 401
rect 812 397 860 402
rect 880 411 1245 413
rect 880 405 885 411
rect 917 405 922 411
rect 926 405 931 411
rect 1005 400 1009 411
rect 753 387 763 391
rect 836 390 841 397
rect 676 377 681 386
rect 759 383 763 387
rect 722 380 763 383
rect 722 377 725 380
rect 759 377 763 380
rect 848 390 853 397
rect 898 390 903 400
rect 961 395 1009 400
rect 1029 409 1154 411
rect 1173 409 1245 411
rect 1390 409 1476 414
rect 1693 509 1701 523
rect 1692 504 1702 509
rect 1029 403 1034 409
rect 1066 403 1071 409
rect 1075 403 1080 409
rect 1149 400 1153 409
rect 898 386 908 390
rect 985 388 990 395
rect 668 373 681 377
rect 693 373 725 377
rect 676 369 681 373
rect 733 372 735 375
rect 665 360 672 361
rect 691 360 696 364
rect 733 361 736 372
rect 750 369 753 372
rect 777 361 780 375
rect 821 376 826 385
rect 904 382 908 386
rect 867 379 908 382
rect 867 376 870 379
rect 904 376 908 379
rect 997 388 1002 395
rect 1047 388 1052 398
rect 1105 395 1153 400
rect 1173 403 1178 409
rect 1210 403 1215 409
rect 1219 403 1224 409
rect 1397 402 1402 409
rect 1129 388 1134 395
rect 1047 384 1057 388
rect 809 373 826 376
rect 818 372 826 373
rect 838 372 870 376
rect 821 368 826 372
rect 878 371 880 374
rect 970 374 975 383
rect 1053 380 1057 384
rect 1016 377 1057 380
rect 1016 374 1019 377
rect 1053 374 1057 377
rect 1141 388 1146 395
rect 1191 388 1196 398
rect 1409 402 1414 409
rect 1447 402 1452 409
rect 1191 384 1201 388
rect 665 355 701 360
rect 665 328 672 355
rect 733 356 780 361
rect 836 359 841 363
rect 878 360 881 371
rect 895 368 898 371
rect 922 360 925 374
rect 952 369 975 374
rect 987 370 1019 374
rect 970 366 975 369
rect 1027 369 1029 372
rect 811 354 846 359
rect 742 346 747 347
rect 765 345 770 347
rect 811 328 818 354
rect 878 355 925 360
rect 985 357 990 361
rect 1027 358 1030 369
rect 1044 366 1047 369
rect 1071 358 1074 372
rect 1114 374 1119 383
rect 1197 380 1201 384
rect 1410 384 1412 388
rect 1410 383 1411 384
rect 1424 380 1429 397
rect 1462 388 1467 397
rect 1447 384 1450 388
rect 1462 383 1465 388
rect 1462 380 1467 383
rect 1160 377 1201 380
rect 1160 374 1163 377
rect 1197 374 1201 377
rect 1095 370 1119 374
rect 1131 370 1163 374
rect 1114 366 1119 370
rect 1171 369 1173 372
rect 954 352 995 357
rect 887 345 892 346
rect 910 345 915 346
rect 955 328 962 352
rect 1027 353 1074 358
rect 1129 357 1134 361
rect 1171 358 1174 369
rect 1188 366 1191 369
rect 1215 358 1218 372
rect 1409 371 1414 375
rect 1447 373 1452 375
rect 1434 371 1453 373
rect 1353 370 1479 371
rect 1353 366 1437 370
rect 1450 368 1479 370
rect 1452 366 1479 368
rect 1353 363 1404 366
rect 1104 352 1139 357
rect 1036 343 1041 344
rect 1059 343 1064 344
rect 1103 328 1112 352
rect 1171 353 1218 358
rect 1180 343 1185 344
rect 1203 343 1208 344
rect 1249 335 1318 339
rect 665 327 1112 328
rect 647 322 1112 327
rect 665 321 672 322
rect 955 320 962 322
rect 1103 303 1111 322
rect 1398 303 1404 363
rect 1103 299 1405 303
rect 1319 131 1323 171
rect 1398 161 1404 299
rect 1442 262 1446 361
rect 1488 274 1496 482
rect 1596 448 1627 449
rect 1548 445 1627 448
rect 1548 443 1599 445
rect 1548 437 1553 443
rect 1557 437 1562 443
rect 1594 437 1599 443
rect 1619 434 1623 445
rect 1693 434 1701 504
rect 1935 509 1944 511
rect 1729 504 1944 509
rect 1935 475 1944 504
rect 2076 475 2083 544
rect 2118 542 2125 544
rect 2408 543 2415 544
rect 1935 469 2084 475
rect 2076 467 2083 469
rect 1576 422 1581 432
rect 1617 429 1701 434
rect 1571 418 1581 422
rect 1624 422 1629 429
rect 1571 414 1575 418
rect 1636 422 1641 429
rect 1674 428 1688 429
rect 1571 411 1612 414
rect 1571 408 1575 411
rect 1609 408 1612 411
rect 1651 408 1656 417
rect 1554 392 1557 406
rect 1599 403 1601 406
rect 1609 404 1639 408
rect 1651 404 1668 408
rect 1581 400 1584 403
rect 1598 392 1601 403
rect 1651 400 1656 404
rect 1554 387 1601 392
rect 1636 391 1641 395
rect 1632 386 1662 391
rect 1564 375 1569 378
rect 1586 375 1592 378
rect 1595 344 1626 345
rect 1547 341 1626 344
rect 1547 339 1598 341
rect 1547 333 1552 339
rect 1556 333 1561 339
rect 1593 333 1598 339
rect 1618 330 1622 341
rect 1693 330 1701 429
rect 1575 318 1580 328
rect 1618 325 1701 330
rect 1570 314 1580 318
rect 1625 318 1630 325
rect 1570 310 1574 314
rect 1637 318 1642 325
rect 1570 307 1611 310
rect 1570 304 1574 307
rect 1608 304 1611 307
rect 1652 304 1657 313
rect 1553 288 1556 302
rect 1598 299 1600 302
rect 1608 300 1640 304
rect 1652 300 1670 304
rect 1580 296 1583 299
rect 1597 288 1600 299
rect 1652 296 1657 300
rect 1553 283 1600 288
rect 1637 287 1642 291
rect 1631 282 1658 287
rect 1488 269 1568 274
rect 1586 262 1591 274
rect 1442 256 1591 262
rect 1533 179 1537 256
rect 1595 248 1626 249
rect 1547 245 1626 248
rect 1547 243 1598 245
rect 1547 237 1552 243
rect 1556 237 1561 243
rect 1593 237 1598 243
rect 1618 234 1622 245
rect 1693 234 1701 325
rect 1575 222 1580 232
rect 1616 229 1701 234
rect 1570 218 1580 222
rect 1624 222 1629 229
rect 1570 214 1574 218
rect 1636 222 1641 229
rect 1570 211 1611 214
rect 1570 208 1574 211
rect 1608 208 1611 211
rect 1651 208 1656 217
rect 1553 192 1556 206
rect 1598 203 1600 206
rect 1608 204 1639 208
rect 1651 204 1805 208
rect 1580 200 1583 203
rect 1597 192 1600 203
rect 1651 200 1656 204
rect 1553 187 1600 192
rect 1636 191 1641 195
rect 1657 191 1665 192
rect 1632 186 1665 191
rect 1657 185 1665 186
rect 1533 178 1563 179
rect 1533 175 1568 178
rect 1659 161 1665 185
rect 1398 156 1665 161
rect 1319 126 1831 131
rect 476 23 641 29
rect 673 6 682 92
rect 299 0 682 6
<< m2contact >>
rect 944 1020 949 1025
rect 895 1010 902 1017
rect 936 995 941 1002
rect 859 984 869 989
rect 944 984 950 989
rect 943 960 949 966
rect 882 929 889 936
rect 669 893 674 900
rect 866 897 872 906
rect 700 891 707 897
rect 795 880 800 886
rect 132 802 141 813
rect 655 864 661 869
rect 795 864 802 869
rect 1071 853 1086 862
rect 655 844 662 849
rect 795 844 802 849
rect 931 846 936 851
rect 186 777 199 787
rect 75 763 86 773
rect 461 761 475 771
rect 186 733 193 739
rect 229 708 234 713
rect 356 733 361 738
rect 227 690 232 695
rect 287 707 294 712
rect 250 690 255 695
rect 304 667 309 672
rect 383 695 390 702
rect 398 693 403 700
rect 458 690 463 695
rect 530 749 538 757
rect 604 823 615 830
rect 655 823 663 829
rect 736 824 750 829
rect 795 826 802 831
rect 578 701 587 715
rect 931 825 937 830
rect 840 789 853 805
rect 655 779 664 786
rect 681 777 690 785
rect 796 782 801 788
rect 899 789 909 798
rect 1077 792 1088 803
rect 1176 786 1187 795
rect 2071 807 2083 818
rect 796 758 801 765
rect 615 743 622 748
rect 961 742 967 750
rect 1116 725 1126 731
rect 1206 717 1211 722
rect 1157 707 1164 714
rect 690 696 695 702
rect 706 696 711 702
rect 754 696 759 703
rect 472 665 477 670
rect 720 666 730 674
rect 755 672 765 680
rect 545 648 561 660
rect 503 599 517 608
rect 224 539 229 544
rect 183 510 190 516
rect 226 486 231 491
rect 353 511 358 516
rect 224 468 229 473
rect 286 482 292 488
rect 247 468 252 473
rect 379 473 388 478
rect 301 445 306 450
rect 455 468 460 473
rect 469 443 474 448
rect 568 647 585 658
rect 548 598 560 610
rect 621 623 633 634
rect 570 581 581 596
rect 541 558 552 569
rect 739 642 751 658
rect 914 629 925 638
rect 1198 692 1203 699
rect 1221 692 1226 699
rect 1012 623 1024 630
rect 1039 623 1051 630
rect 779 579 789 586
rect 815 577 828 587
rect 716 562 727 573
rect 958 560 970 574
rect 1102 568 1117 577
rect 1318 554 1326 561
rect 573 531 585 541
rect 651 532 662 541
rect 1663 762 1676 775
rect 1991 763 1998 771
rect 2618 794 2628 803
rect 2186 778 2194 785
rect 2114 770 2124 777
rect 2132 758 2142 766
rect 2262 774 2271 780
rect 2766 771 2776 781
rect 2281 759 2289 765
rect 1887 691 1892 696
rect 1980 698 1986 705
rect 1934 681 1941 688
rect 2023 691 2028 696
rect 2118 699 2124 706
rect 1872 666 1877 673
rect 1895 666 1900 673
rect 2070 681 2077 688
rect 2169 693 2174 698
rect 2264 700 2270 707
rect 2216 683 2223 690
rect 2316 693 2321 698
rect 2420 700 2427 708
rect 2008 666 2013 673
rect 2031 666 2036 673
rect 2154 668 2159 675
rect 2177 668 2182 675
rect 2363 683 2370 690
rect 2528 692 2533 697
rect 2281 667 2289 673
rect 2301 668 2306 675
rect 2324 668 2329 675
rect 2575 682 2582 689
rect 2664 692 2669 697
rect 2513 667 2518 674
rect 2536 667 2541 674
rect 2711 682 2718 689
rect 2810 694 2815 699
rect 2857 684 2864 691
rect 2957 694 2962 699
rect 2649 667 2654 674
rect 2672 667 2677 674
rect 2795 669 2800 676
rect 2818 669 2823 676
rect 3004 684 3011 691
rect 2942 669 2947 676
rect 2965 669 2970 676
rect 1887 583 1892 588
rect 1993 591 1998 597
rect 1934 573 1941 580
rect 2031 583 2036 588
rect 2133 589 2139 596
rect 1832 553 1838 560
rect 1872 557 1877 565
rect 1895 558 1900 565
rect 660 480 667 486
rect 759 471 764 476
rect 815 481 821 486
rect 710 461 717 468
rect 906 471 911 476
rect 959 478 966 484
rect 153 400 160 407
rect 198 401 205 408
rect 480 360 489 370
rect 144 348 152 354
rect 45 300 50 305
rect 161 326 168 332
rect 356 326 361 331
rect 228 299 233 305
rect 227 283 232 288
rect 147 267 153 273
rect 186 267 192 272
rect 226 255 231 261
rect 143 243 151 249
rect 288 298 293 303
rect 250 283 255 288
rect 304 260 309 265
rect 383 288 391 293
rect 458 283 463 288
rect 472 258 477 263
rect 542 432 554 443
rect 572 438 583 448
rect 751 446 756 453
rect 774 446 779 453
rect 857 461 864 468
rect 1052 469 1057 474
rect 1103 476 1109 481
rect 898 446 903 453
rect 1003 459 1010 466
rect 1188 469 1193 474
rect 921 446 926 453
rect 1044 444 1049 451
rect 1067 444 1072 451
rect 1139 459 1146 466
rect 1180 444 1185 451
rect 1203 444 1208 451
rect 541 376 551 389
rect 535 349 545 357
rect 635 373 641 378
rect 620 324 630 334
rect 501 225 510 232
rect 502 196 509 203
rect 510 168 516 176
rect 186 151 193 157
rect 356 151 361 156
rect 228 125 233 130
rect 227 108 232 113
rect 288 123 294 128
rect 250 108 255 113
rect 378 113 388 118
rect 304 85 309 90
rect 458 108 463 113
rect 472 83 477 88
rect 617 95 626 107
rect 476 38 485 48
rect 1580 513 1585 518
rect 1660 522 1666 527
rect 2078 573 2085 580
rect 2180 585 2185 590
rect 2282 592 2288 598
rect 2227 575 2234 582
rect 2325 586 2330 591
rect 2407 592 2415 599
rect 2372 576 2379 583
rect 2016 558 2021 565
rect 2039 558 2044 565
rect 2165 560 2170 567
rect 2188 560 2193 567
rect 2310 560 2315 567
rect 2333 561 2338 568
rect 1627 504 1634 510
rect 1488 482 1496 490
rect 1565 489 1570 496
rect 1656 501 1665 510
rect 1832 518 1838 523
rect 1588 490 1593 496
rect 662 371 668 377
rect 750 364 755 369
rect 804 373 809 378
rect 701 354 708 361
rect 895 363 900 368
rect 945 369 952 374
rect 742 339 747 346
rect 765 338 770 345
rect 846 353 853 360
rect 1044 361 1049 366
rect 1090 370 1095 375
rect 1405 383 1410 388
rect 1429 383 1435 388
rect 1442 383 1447 388
rect 1465 383 1473 388
rect 887 338 892 345
rect 910 338 915 345
rect 995 351 1002 358
rect 1188 361 1193 366
rect 1337 363 1353 375
rect 1036 336 1041 343
rect 1059 336 1064 343
rect 1139 351 1146 358
rect 1180 336 1185 343
rect 1203 335 1208 343
rect 1244 335 1249 341
rect 1318 335 1323 341
rect 1441 361 1447 366
rect 1319 171 1326 177
rect 1720 503 1729 512
rect 1579 395 1584 400
rect 1624 386 1632 391
rect 1564 370 1569 375
rect 1586 369 1592 375
rect 1670 300 1678 306
rect 1578 291 1583 296
rect 1623 282 1631 288
rect 1578 195 1583 200
rect 1805 203 1815 210
rect 1624 185 1632 191
rect 1586 171 1591 178
rect 1831 123 1839 136
rect 671 92 685 107
rect 288 0 299 11
<< metal2 >>
rect 918 1020 944 1023
rect 918 1016 923 1020
rect 902 1011 923 1016
rect 632 995 936 998
rect 632 993 941 995
rect 633 914 636 993
rect 869 984 888 989
rect 883 936 888 984
rect 944 966 947 984
rect 46 911 636 914
rect 46 761 50 911
rect 655 893 669 895
rect 872 899 906 904
rect 655 891 674 893
rect 707 892 824 895
rect 754 891 824 892
rect 655 869 659 891
rect 796 869 800 880
rect 342 856 1071 860
rect 125 804 132 809
rect 343 788 348 856
rect 554 825 604 829
rect 655 829 660 844
rect 742 829 746 856
rect 796 831 800 844
rect 931 830 935 846
rect 1925 843 1932 844
rect 1925 842 2193 843
rect 1925 838 2194 842
rect 571 815 1257 819
rect 199 777 283 785
rect 178 769 234 770
rect 86 767 234 769
rect 343 767 349 788
rect 86 764 349 767
rect 86 763 184 764
rect 45 680 50 761
rect 45 305 49 680
rect 154 407 158 740
rect 186 516 189 733
rect 229 713 234 764
rect 364 761 461 767
rect 364 758 471 761
rect 364 738 369 758
rect 361 733 383 738
rect 232 690 250 695
rect 288 590 293 707
rect 377 695 383 733
rect 390 695 398 700
rect 458 695 463 758
rect 571 754 580 815
rect 731 798 840 799
rect 645 793 840 798
rect 645 792 759 793
rect 538 749 580 754
rect 615 779 655 784
rect 681 785 688 792
rect 853 793 856 799
rect 1008 794 1077 797
rect 909 792 1077 794
rect 909 789 1081 792
rect 615 748 621 779
rect 796 765 800 782
rect 961 750 966 778
rect 1116 731 1120 792
rect 1177 720 1182 786
rect 1251 774 1257 815
rect 1925 809 1932 838
rect 1612 803 1932 809
rect 1955 817 1960 818
rect 1955 811 2071 817
rect 1177 717 1206 720
rect 556 706 578 712
rect 304 625 309 667
rect 462 665 472 669
rect 462 625 468 665
rect 556 660 562 706
rect 1177 713 1185 717
rect 1164 708 1185 713
rect 1250 697 1257 774
rect 1226 694 1257 697
rect 1226 693 1254 694
rect 1198 688 1203 692
rect 714 666 720 672
rect 561 648 562 660
rect 585 647 739 655
rect 304 624 610 625
rect 304 620 612 624
rect 633 629 720 630
rect 633 623 721 629
rect 457 619 612 620
rect 596 617 612 619
rect 517 599 548 606
rect 288 585 570 590
rect 186 359 189 510
rect 226 491 229 539
rect 361 536 468 545
rect 361 516 366 536
rect 358 511 380 516
rect 229 468 247 473
rect 205 402 232 406
rect 161 355 189 359
rect 161 354 164 355
rect 152 348 164 354
rect 228 352 232 402
rect 287 383 291 482
rect 374 478 380 511
rect 374 473 379 478
rect 455 473 460 536
rect 301 403 306 445
rect 459 443 469 447
rect 542 443 548 558
rect 575 448 580 531
rect 459 403 465 443
rect 301 400 465 403
rect 301 398 565 400
rect 454 397 565 398
rect 287 379 541 383
rect 398 364 480 368
rect 161 332 164 348
rect 200 349 232 352
rect 200 337 205 349
rect 186 334 205 337
rect 146 267 147 272
rect 146 249 149 267
rect 161 249 164 326
rect 186 272 190 334
rect 228 305 232 349
rect 364 351 471 360
rect 364 331 369 351
rect 361 326 383 331
rect 232 283 250 288
rect 161 245 189 249
rect 186 157 189 245
rect 228 130 231 255
rect 289 200 293 298
rect 377 288 383 326
rect 458 288 463 351
rect 304 218 309 260
rect 462 258 472 262
rect 462 218 468 258
rect 537 230 542 349
rect 560 328 565 397
rect 510 227 542 230
rect 510 226 541 227
rect 304 216 468 218
rect 558 217 565 328
rect 600 290 610 617
rect 634 591 640 592
rect 634 586 706 591
rect 634 488 640 586
rect 699 557 705 586
rect 716 573 721 623
rect 758 557 763 672
rect 1613 662 1621 803
rect 1955 789 1960 811
rect 2188 816 2194 838
rect 802 652 1621 662
rect 781 563 787 579
rect 699 553 763 557
rect 780 539 787 563
rect 662 532 787 539
rect 620 487 656 488
rect 620 486 664 487
rect 620 482 660 486
rect 620 334 628 482
rect 633 481 660 482
rect 733 471 759 474
rect 733 467 738 471
rect 717 462 738 467
rect 803 451 810 652
rect 1613 651 1621 652
rect 1635 781 1960 789
rect 1979 785 2156 790
rect 2188 785 2193 816
rect 2628 794 2629 803
rect 2246 785 2456 790
rect 1979 784 2006 785
rect 1635 641 1641 781
rect 943 634 1642 641
rect 815 555 819 577
rect 918 555 923 629
rect 815 551 924 555
rect 815 486 819 551
rect 880 471 906 474
rect 880 467 885 471
rect 864 462 885 467
rect 779 448 810 451
rect 779 447 807 448
rect 751 428 756 446
rect 898 428 903 446
rect 943 450 950 634
rect 1007 623 1012 629
rect 1024 623 1039 630
rect 959 554 963 560
rect 1007 554 1014 623
rect 1664 612 1670 762
rect 1980 705 1986 784
rect 2118 777 2123 778
rect 1892 691 1918 694
rect 1913 687 1918 691
rect 1913 682 1934 687
rect 1092 604 1670 612
rect 1772 661 1777 663
rect 1872 662 1877 666
rect 1855 661 1877 662
rect 1772 657 1877 661
rect 1772 656 1861 657
rect 959 548 1015 554
rect 959 484 963 548
rect 1026 469 1052 472
rect 1026 465 1031 469
rect 1010 460 1031 465
rect 926 446 950 450
rect 921 445 948 446
rect 1092 447 1097 604
rect 1253 590 1260 591
rect 1772 590 1777 656
rect 1895 650 1900 666
rect 1991 670 1996 763
rect 2118 706 2123 770
rect 2151 758 2156 785
rect 2246 758 2250 785
rect 2028 691 2054 694
rect 2049 687 2054 691
rect 2049 682 2070 687
rect 1991 666 2008 670
rect 2134 671 2139 758
rect 2151 754 2250 758
rect 2264 707 2269 774
rect 2174 693 2200 696
rect 2195 689 2200 693
rect 2195 684 2216 689
rect 2134 668 2154 671
rect 2134 667 2159 668
rect 2139 666 2155 667
rect 1991 665 2005 666
rect 1991 664 1996 665
rect 2031 650 2036 666
rect 2177 650 2182 668
rect 2281 673 2285 759
rect 2421 708 2427 755
rect 2321 693 2347 696
rect 2342 689 2347 693
rect 2342 684 2363 689
rect 2289 671 2297 672
rect 2289 668 2301 671
rect 2289 667 2306 668
rect 2324 650 2329 668
rect 2450 662 2456 785
rect 2533 692 2559 695
rect 2554 688 2559 692
rect 2554 683 2575 688
rect 2513 662 2518 667
rect 2450 657 2518 662
rect 2625 671 2629 794
rect 2776 771 2777 780
rect 2669 692 2695 695
rect 2690 688 2695 692
rect 2690 683 2711 688
rect 2624 667 2649 671
rect 2771 673 2777 771
rect 2915 753 2916 760
rect 2815 694 2841 697
rect 2836 690 2841 694
rect 2836 685 2857 690
rect 2771 672 2789 673
rect 2771 669 2795 672
rect 2771 668 2800 669
rect 2911 672 2916 753
rect 2962 694 2988 697
rect 2983 690 2988 694
rect 2983 685 3004 690
rect 1253 584 1777 590
rect 1103 563 1109 568
rect 1103 557 1199 563
rect 1103 481 1109 557
rect 1162 469 1188 472
rect 1162 465 1167 469
rect 1146 460 1167 465
rect 1072 444 1098 447
rect 1044 428 1049 444
rect 1180 428 1185 444
rect 1253 446 1260 584
rect 1772 582 1777 584
rect 1810 647 2329 650
rect 1208 444 1260 446
rect 1203 441 1260 444
rect 1318 500 1323 554
rect 1810 536 1814 647
rect 1892 583 1918 586
rect 1913 579 1918 583
rect 1993 580 1998 591
rect 2415 594 2456 599
rect 2036 583 2062 586
rect 1913 574 1934 579
rect 2057 579 2062 583
rect 2057 574 2078 579
rect 2133 568 2139 589
rect 2185 585 2211 588
rect 2206 581 2211 585
rect 2206 576 2227 581
rect 2284 570 2288 592
rect 2330 586 2356 589
rect 2351 582 2356 586
rect 2351 577 2372 582
rect 1861 560 1872 561
rect 1838 557 1872 560
rect 1895 536 1900 558
rect 2010 558 2016 561
rect 2010 557 2021 558
rect 2039 536 2044 558
rect 2159 560 2165 563
rect 2159 559 2170 560
rect 2188 536 2193 560
rect 2306 560 2310 564
rect 2333 536 2338 561
rect 1810 533 2338 536
rect 1666 523 1683 527
rect 1810 526 1814 533
rect 2333 532 2338 533
rect 1806 523 1814 526
rect 1585 513 1611 516
rect 1606 509 1611 513
rect 1606 505 1627 509
rect 1606 504 1618 505
rect 751 425 1270 428
rect 641 373 662 377
rect 724 364 750 367
rect 804 368 807 373
rect 724 360 729 364
rect 869 363 895 366
rect 708 355 729 360
rect 869 359 874 363
rect 853 354 874 359
rect 945 361 948 369
rect 1018 361 1044 364
rect 1018 357 1023 361
rect 1002 352 1023 357
rect 1090 350 1094 370
rect 1162 361 1188 364
rect 1162 357 1167 361
rect 1146 352 1167 357
rect 742 314 747 339
rect 770 339 792 343
rect 887 314 892 338
rect 915 338 931 340
rect 910 336 931 338
rect 1064 336 1074 340
rect 1036 314 1041 336
rect 1180 314 1185 336
rect 1208 335 1244 339
rect 1266 314 1270 425
rect 1318 371 1324 500
rect 1433 482 1488 487
rect 1565 487 1570 489
rect 1496 482 1570 487
rect 1433 390 1438 482
rect 1588 472 1593 490
rect 1520 465 1593 472
rect 1433 388 1437 390
rect 1520 388 1527 465
rect 1584 395 1607 398
rect 1388 383 1405 388
rect 1435 383 1437 388
rect 1473 383 1527 388
rect 1602 391 1607 395
rect 1611 391 1616 504
rect 1665 504 1720 510
rect 1602 386 1624 391
rect 1318 364 1337 371
rect 1388 357 1394 383
rect 1442 366 1446 383
rect 1520 371 1527 383
rect 1520 370 1564 371
rect 1520 364 1569 370
rect 1586 357 1592 369
rect 1388 353 1592 357
rect 1388 352 1394 353
rect 742 311 1270 314
rect 742 310 747 311
rect 600 287 1090 290
rect 600 286 610 287
rect 896 266 900 271
rect 895 263 946 266
rect 953 263 954 266
rect 895 262 954 263
rect 772 248 805 251
rect 772 247 810 248
rect 558 216 616 217
rect 896 216 900 262
rect 1080 232 1247 238
rect 304 213 551 216
rect 289 196 502 200
rect 364 176 471 185
rect 510 176 516 182
rect 364 156 369 176
rect 361 151 383 156
rect 232 108 250 113
rect 288 28 292 123
rect 377 118 383 151
rect 377 113 378 118
rect 458 113 463 176
rect 304 43 309 85
rect 462 83 472 87
rect 462 44 468 83
rect 461 43 476 44
rect 304 38 476 43
rect 542 42 551 213
rect 558 213 903 216
rect 558 210 616 213
rect 940 216 1218 218
rect 940 212 1219 216
rect 800 184 1182 188
rect 626 95 671 104
rect 749 44 759 45
rect 631 43 759 44
rect 571 42 759 43
rect 542 39 759 42
rect 542 38 749 39
rect 1177 48 1182 184
rect 1209 81 1219 212
rect 1242 211 1247 232
rect 1242 133 1248 211
rect 1266 150 1270 311
rect 1319 177 1322 335
rect 1428 171 1432 353
rect 1583 291 1607 294
rect 1602 287 1607 291
rect 1611 287 1616 386
rect 1669 300 1670 304
rect 1678 300 1719 304
rect 1602 282 1623 287
rect 1583 195 1606 198
rect 1602 191 1606 195
rect 1611 191 1616 282
rect 1602 186 1624 191
rect 1428 168 1591 171
rect 1586 167 1591 168
rect 1713 150 1719 300
rect 1806 210 1810 523
rect 2154 522 2158 523
rect 1834 495 1837 518
rect 1266 145 1719 150
rect 1713 144 1719 145
rect 1833 136 1837 495
rect 2006 458 2010 493
rect 2154 468 2158 516
rect 2364 471 2367 526
rect 2536 490 2541 667
rect 2672 505 2677 667
rect 2818 521 2823 669
rect 2910 669 2942 672
rect 2910 668 2947 669
rect 2965 651 2970 669
rect 2966 602 2970 651
rect 1892 449 2010 458
rect 2153 459 2158 468
rect 2177 466 2367 471
rect 1243 105 1248 133
rect 1892 105 1897 449
rect 1919 419 1928 421
rect 2153 419 2157 459
rect 1919 411 2160 419
rect 1243 99 1902 105
rect 1209 76 1218 81
rect 1919 76 1928 411
rect 2177 397 2189 466
rect 1966 385 2189 397
rect 1209 66 1930 76
rect 1919 64 1928 66
rect 1967 48 1977 385
rect 1177 39 1977 48
rect 288 11 293 28
<< m3contact >>
rect 906 898 913 904
rect 824 888 837 896
rect 113 801 125 813
rect 546 824 554 833
rect 283 776 299 788
rect 152 740 160 748
rect 631 790 645 801
rect 1114 792 1127 799
rect 959 778 967 783
rect 1197 682 1205 688
rect 706 666 714 674
rect 387 364 398 372
rect 2421 755 2429 763
rect 2906 753 2915 763
rect 1199 557 1207 563
rect 2456 592 2466 600
rect 1993 574 1998 580
rect 2004 555 2010 563
rect 2132 561 2139 568
rect 2153 556 2159 564
rect 2283 563 2289 570
rect 2298 558 2306 568
rect 2361 526 2368 532
rect 804 363 809 368
rect 945 356 950 361
rect 1090 345 1095 350
rect 792 339 797 345
rect 931 335 938 341
rect 1074 336 1080 343
rect 1090 286 1095 291
rect 946 263 953 269
rect 763 246 772 254
rect 805 248 812 254
rect 1072 232 1080 242
rect 510 182 517 190
rect 931 212 940 221
rect 795 184 800 192
rect 759 36 771 49
rect 2153 516 2160 522
rect 2004 493 2012 500
rect 2965 593 2975 602
rect 2816 513 2826 521
rect 2669 498 2679 505
rect 2536 482 2543 490
<< metal3 >>
rect 913 898 1033 903
rect 1029 889 1033 898
rect 829 886 1000 888
rect 1029 886 1119 889
rect 829 884 1001 886
rect 1029 884 1121 886
rect 154 831 157 832
rect 152 826 546 831
rect 116 393 120 801
rect 154 748 157 826
rect 390 797 394 799
rect 535 797 631 798
rect 389 793 631 797
rect 390 785 394 793
rect 535 791 631 793
rect 299 776 395 785
rect 997 783 1001 884
rect 1116 799 1121 884
rect 967 778 1002 783
rect 2429 761 2439 762
rect 2429 756 2906 761
rect 2429 755 2439 756
rect 607 601 615 603
rect 707 601 712 666
rect 606 594 713 601
rect 580 410 587 412
rect 607 410 615 594
rect 1199 563 1202 682
rect 2461 600 2965 602
rect 2466 593 2965 600
rect 1993 485 1998 574
rect 2005 500 2010 555
rect 2132 505 2139 561
rect 2154 522 2158 556
rect 2283 518 2289 563
rect 2300 530 2303 558
rect 2300 527 2361 530
rect 2283 513 2816 518
rect 2132 499 2669 505
rect 1993 482 2536 485
rect 1993 481 2542 482
rect 580 403 616 410
rect 116 389 248 393
rect 240 369 245 389
rect 240 365 387 369
rect 580 292 587 403
rect 797 339 798 344
rect 579 188 587 292
rect 517 182 587 188
rect 761 246 763 252
rect 761 49 766 246
rect 795 192 798 339
rect 806 254 809 363
rect 931 221 937 335
rect 946 269 949 356
rect 1073 336 1074 338
rect 1073 242 1079 336
rect 1090 291 1094 345
<< labels >>
rlabel metal1 1426 386 1426 386 1 S0c
rlabel metal1 1411 386 1411 386 1 S0
rlabel metal1 1449 387 1449 387 1 S1
rlabel metal1 1665 406 1665 406 1 D1
rlabel metal1 1659 525 1659 525 1 D0
rlabel metal1 1667 206 1667 206 1 D3
rlabel metal1 1576 189 1576 189 1 DEC_AND_NODE_4
rlabel metal1 1576 212 1576 212 1 DEC_D3_NAND
rlabel metal1 1668 302 1668 302 1 D2
rlabel metal1 1577 285 1577 285 1 DEC_AND_NODE_3
rlabel metal1 1577 308 1577 308 1 DEC_D2_NAND
rlabel metal1 1579 389 1579 389 1 Dec_AND_node_2
rlabel metal1 1580 412 1580 412 1 DEC_D1_NAND
rlabel metal1 1575 531 1575 531 1 DEC_D0_NAND
rlabel metal1 1580 508 1580 508 1 Dec_AND_node_1
rlabel m2contact 1468 386 1468 386 1 S1c
rlabel metal1 1468 368 1468 368 1 gnd
rlabel metal1 1444 412 1444 412 1 vdd
rlabel metal2 1867 559 1867 559 1 B3
rlabel m3contact 2008 560 2008 560 1 B2
rlabel metal2 2160 562 2160 562 1 B1
rlabel metal1 2326 580 2326 580 1 ander_node_5
rlabel metal1 2178 580 2178 580 1 ander_node_6
rlabel metal1 2029 576 2029 576 1 ander_node_7
rlabel metal1 1884 578 1884 578 1 ander_node_8
rlabel metal1 2360 597 2360 597 1 and_b0e_nand
rlabel metal1 2225 596 2225 596 1 and_b1e_nand
rlabel metal1 2071 593 2071 593 1 and_b2e_nand
rlabel metal1 1923 593 1923 593 1 and_b3e_nand
rlabel metal1 2404 597 2404 597 1 and_b0e
rlabel metal1 2260 596 2260 596 1 and_b1e
rlabel metal1 2112 593 2112 593 1 and_b2e
rlabel metal1 1968 594 1968 594 1 and_b3e
rlabel metal1 2395 703 2395 703 1 and_a0e
rlabel metal1 2248 703 2248 703 1 and_a1e
rlabel metal1 2101 701 2101 701 1 and_a2e
rlabel metal1 1966 702 1966 702 1 and_a3e
rlabel metal1 2358 703 2358 703 1 and_a0e_nand
rlabel metal1 2212 704 2212 704 1 and_a1e_nand
rlabel metal1 2069 702 2069 702 1 and_a2e_nand
rlabel metal1 1925 703 1925 703 1 and_a3e_nand
rlabel metal1 2315 687 2315 687 1 ander_node_4
rlabel metal1 2168 687 2168 687 1 ander_node_3
rlabel metal1 2022 686 2022 686 1 ander_node_2
rlabel metal1 1886 685 1886 685 1 ander_node_1
rlabel metal2 2295 669 2295 669 1 A0
rlabel metal2 2149 669 2149 669 1 A1
rlabel metal2 2002 667 2002 667 1 A2
rlabel metal2 1874 662 1874 662 1 A3
rlabel metal1 2526 687 2526 687 1 ander_node_9
rlabel metal1 2660 687 2660 687 1 ander_node_10
rlabel metal1 2810 690 2810 690 1 ander_node_11
rlabel metal1 2954 687 2954 687 1 ander_node_12
rlabel metal1 2567 703 2567 703 1 A3_and_B3_nand
rlabel metal1 2695 704 2695 704 1 A2_and_B2_nand
rlabel metal1 2850 705 2850 705 1 A1_and_B1_nand
rlabel metal1 2990 705 2990 705 1 A0_and_B0_nand
rlabel metal1 2608 703 2608 703 1 A3_and_B3
rlabel metal1 2744 703 2744 703 1 A2_and_B2
rlabel metal1 2889 705 2889 705 1 A1_and_B1
rlabel metal1 3037 705 3037 705 1 A0_and_B0
rlabel metal1 1197 464 1197 464 1 compare_node_1
rlabel metal1 1058 464 1058 464 1 compare_node_2
rlabel metal1 912 465 912 465 1 compare_node_3
rlabel metal1 766 465 766 465 1 compare_node_4
rlabel metal1 757 359 757 359 1 compare_node_5
rlabel metal1 901 357 901 357 1 compare_node_6
rlabel metal1 1051 354 1051 354 1 compare_node_7
rlabel metal1 1194 354 1194 354 1 compare_node_8
rlabel metal1 1197 495 1197 495 1 compare_A3e_nand
rlabel metal1 1063 494 1063 494 1 compare_A2e_nand
rlabel metal1 917 493 917 493 1 compare_A1e_nand
rlabel metal1 769 497 769 497 1 compare_A0e_nand
rlabel metal1 761 390 761 390 1 compare_B0e_nand
rlabel metal1 906 387 906 387 1 compare_B1e_nand
rlabel metal1 1054 386 1054 386 1 compare_B2e_nand
rlabel metal1 1199 386 1199 386 1 compare_B3e_nand
rlabel metal1 1113 480 1113 480 1 compare_A3e
rlabel metal1 978 481 978 481 1 compare_A2e
rlabel metal1 834 481 834 481 1 compare_A1e
rlabel metal1 685 483 685 483 1 compare_A0e
rlabel metal1 677 375 677 375 1 compare_B0e
rlabel metal1 823 374 823 374 1 compare_B1e
rlabel metal1 972 371 972 371 1 compare_B2e
rlabel metal1 1117 372 1117 372 1 compare_B3e
rlabel pdiffusion 335 720 335 720 1 xnor_1
rlabel ndiffusion 335 680 335 680 1 xnor_2
rlabel metal1 396 709 396 709 1 xor_1
rlabel ndiffusion 417 720 417 720 1 xnor_3
rlabel pdiffusion 417 680 417 680 1 xnor_4
rlabel metal1 425 634 425 634 1 A3c
rlabel metal1 382 751 382 751 1 B3c
rlabel pdiffusion 330 498 330 498 1 xnor_5
rlabel ndiffusion 333 458 333 458 1 xnor_6
rlabel ndiffusion 416 498 416 498 1 xnor_7
rlabel pdiffusion 412 457 412 457 1 xnor_8
rlabel metal1 424 409 424 409 1 A2c
rlabel metal1 383 531 383 531 1 B2c
rlabel metal1 383 346 383 346 1 B1c
rlabel metal1 417 223 417 223 1 A1c
rlabel pdiffusion 335 312 335 312 1 xnor_9
rlabel ndiffusion 338 273 338 273 1 xnor_10
rlabel pdiffusion 416 273 416 273 1 xnor_11
rlabel ndiffusion 418 313 418 313 1 xnor_12
rlabel metal1 385 485 385 485 1 xor_2
rlabel metal1 390 301 390 301 1 xor_3
rlabel metal1 393 170 393 170 1 B0c
rlabel metal1 417 49 417 49 1 A0c
rlabel metal1 393 127 393 127 1 xor_4
rlabel pdiffusion 334 138 334 138 1 xnor_13
rlabel ndiffusion 336 97 336 97 1 xnor_14
rlabel ndiffusion 418 137 418 137 1 xnor_15
rlabel pdiffusion 418 98 418 98 1 xnor_16
rlabel ndiffusion 88 290 88 290 1 A_compare_B_node_3
rlabel ndiffusion 105 291 105 291 1 A_compare_B_node_2
rlabel ndiffusion 120 291 120 291 1 A_compare_B_node_1
rlabel metal1 5 315 5 315 3 A_equal_B
rlabel metal1 51 303 51 303 1 A_equal_B_c
rlabel metal1 94 373 94 373 1 A2e_xnor_B2e
rlabel metal1 223 711 223 711 1 A3e_xnor_B3e
rlabel metal1 222 303 222 303 1 A1e_xnor_B1e
rlabel metal1 223 127 223 127 1 A0e_xnor_B0e
rlabel metal2 2307 561 2307 561 1 B0
rlabel metal1 1214 712 1214 712 1 A_greater_B_node_1
rlabel metal1 1126 728 1126 728 1 A3_and_B3c
rlabel metal1 1211 744 1211 744 1 A3_nand_B3c
rlabel ndiffusion 1070 720 1070 720 1 A_greater_B_node_2
rlabel ndiffusion 1054 720 1054 720 1 A_greater_B_node_3
rlabel metal1 1024 728 1024 728 1 A3_eq_B3_A2_gt_B2_c
rlabel metal1 969 746 969 746 1 A3_eq_B3_A2_gt_B2
rlabel ndiffusion 928 721 928 721 1 A_greater_B_node_5
rlabel ndiffusion 907 722 907 722 1 A_greater_B_node_6
rlabel ndiffusion 891 720 891 720 1 A_greater_B_node_7
rlabel metal1 866 734 866 734 1 A3_eq_B3_A2_eq_B2_A1_gt_B1_c
rlabel metal1 812 747 812 747 1 A3_eq_B3_A2_eq_B2_A1_gt_B1
rlabel ndiffusion 734 723 734 723 1 A_greater_B_node_9
rlabel ndiffusion 715 722 715 722 1 A_greater_B_node_10
rlabel ndiffusion 699 722 699 722 1 A_greater_B_node_11
rlabel metal1 675 732 675 732 1 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c
rlabel metal1 622 746 622 746 1 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0
rlabel ndiffusion 750 721 750 721 1 A_greater_B_node_8
rlabel pdiffusion 710 959 710 959 1 A_GT_B_node_1
rlabel pdiffusion 694 958 694 958 1 A_GT_B_node_2
rlabel pdiffusion 677 960 677 960 1 A_GT_B_node_3
rlabel metal1 750 933 750 933 1 A_GT_B_c
rlabel metal1 792 950 792 950 1 A_GT_B
rlabel metal1 948 1014 948 1014 1 A_LS_B_node_1
rlabel metal1 954 1045 954 1045 1 A_LS_B_nand
rlabel metal1 864 1031 864 1031 1 A_LS_B
<< end >>
