magic
tech scmos
timestamp 1701523217
<< nwell >>
rect 863 1035 909 1054
rect 923 1051 984 1068
rect 647 972 731 973
rect 647 953 798 972
rect 809 954 855 973
rect 647 943 752 953
rect 666 769 776 770
rect 855 769 954 770
rect 620 750 776 769
rect 809 750 954 769
rect 967 750 1013 769
rect 674 741 776 750
rect 855 741 954 750
rect 1020 737 1097 769
rect 297 733 361 734
rect 186 714 232 733
rect 257 714 361 733
rect 1125 732 1171 751
rect 1185 748 1246 765
rect 1853 722 1913 739
rect 308 707 361 714
rect 309 706 361 707
rect 1927 706 1973 725
rect 1988 722 2049 739
rect 2063 706 2109 725
rect 2134 724 2195 741
rect 2209 708 2255 727
rect 2282 724 2342 741
rect 2356 708 2402 727
rect 2493 723 2554 740
rect 2568 707 2614 726
rect 2629 723 2690 740
rect 2704 707 2750 726
rect 2775 725 2836 742
rect 2850 709 2896 728
rect 2922 725 2983 742
rect 2997 709 3043 728
rect 376 667 443 695
rect 458 671 504 690
rect 1852 614 1913 631
rect 1927 598 1973 617
rect 1996 614 2057 631
rect 2071 598 2117 617
rect 2145 616 2206 633
rect 2220 600 2266 619
rect 2290 617 2351 634
rect 2365 601 2411 620
rect 1545 544 1606 561
rect 1618 529 1664 548
rect 294 511 358 512
rect 183 492 229 511
rect 254 492 358 511
rect 305 485 358 492
rect 678 486 724 505
rect 738 502 799 519
rect 825 486 871 505
rect 885 502 946 519
rect 306 484 358 485
rect 971 484 1017 503
rect 1031 500 1092 517
rect 1107 484 1153 503
rect 1167 500 1228 517
rect 380 473 403 478
rect 373 445 440 473
rect 455 449 501 468
rect 1544 426 1605 443
rect 2253 434 2314 451
rect 669 379 715 398
rect 729 395 790 412
rect 814 378 860 397
rect 874 394 935 411
rect 1617 410 1663 429
rect 2328 418 2374 437
rect 2389 434 2450 451
rect 2464 418 2510 437
rect 2535 436 2596 453
rect 2610 420 2656 439
rect 2682 436 2743 453
rect 2757 420 2803 439
rect 963 376 1009 395
rect 1023 392 1084 409
rect 1107 376 1153 395
rect 1167 392 1228 409
rect 1390 390 1474 409
rect 2055 375 2101 376
rect 1990 357 2101 375
rect 1990 355 2055 357
rect 49 338 147 339
rect 3 319 147 338
rect 297 326 361 327
rect 49 310 147 319
rect 161 307 232 326
rect 257 307 361 326
rect 1543 322 1604 339
rect 2253 326 2314 343
rect 308 300 361 307
rect 1618 306 1664 325
rect 2328 310 2374 329
rect 2397 326 2458 343
rect 2472 310 2518 329
rect 2546 328 2607 345
rect 2621 312 2667 331
rect 2691 329 2752 346
rect 2766 313 2812 332
rect 309 299 361 300
rect 388 291 406 293
rect 383 288 406 291
rect 376 260 443 288
rect 458 264 504 283
rect 1543 226 1604 243
rect 1616 210 1663 229
rect 297 151 361 152
rect 186 132 232 151
rect 257 132 361 151
rect 308 125 361 132
rect 309 124 361 125
rect 2053 121 2117 122
rect 379 113 406 118
rect 376 85 443 113
rect 458 89 504 108
rect 2009 102 2117 121
rect 2064 95 2117 102
rect 2065 94 2117 95
rect 2147 83 2162 88
rect 2147 74 2199 83
rect 2132 55 2199 74
rect 2214 59 2260 78
rect 1461 -4 1507 15
rect 1514 -14 1598 16
rect 2047 -62 2111 -61
rect 2003 -81 2111 -62
rect 2058 -88 2111 -81
rect 2059 -89 2111 -88
rect 2141 -100 2156 -95
rect 1287 -137 1333 -118
rect 1347 -121 1408 -104
rect 1433 -139 1479 -120
rect 1493 -123 1554 -106
rect 1569 -139 1615 -120
rect 1629 -123 1690 -106
rect 2141 -109 2193 -100
rect 2126 -128 2193 -109
rect 2208 -124 2254 -105
rect 2035 -234 2099 -233
rect 1378 -251 1451 -250
rect 1485 -251 1497 -249
rect 1716 -251 1784 -250
rect 1378 -270 1500 -251
rect 1716 -270 1838 -251
rect 1991 -253 2099 -234
rect 2046 -260 2099 -253
rect 2047 -261 2099 -260
rect 1378 -277 1431 -270
rect 1716 -277 1769 -270
rect 2129 -272 2144 -267
rect 1378 -278 1430 -277
rect 1716 -278 1768 -277
rect 2129 -281 2181 -272
rect 1333 -289 1348 -284
rect 1671 -289 1686 -284
rect 1235 -313 1281 -294
rect 1296 -298 1348 -289
rect 1296 -317 1363 -298
rect 1573 -313 1619 -294
rect 1634 -298 1686 -289
rect 1634 -317 1701 -298
rect 2114 -300 2181 -281
rect 2196 -296 2242 -277
rect 2026 -418 2090 -417
rect 1982 -437 2090 -418
rect 2037 -444 2090 -437
rect 2038 -445 2090 -444
rect 2120 -456 2135 -451
rect 2120 -465 2172 -456
rect 2105 -484 2172 -465
rect 2187 -480 2233 -461
<< ntransistor >>
rect 936 1028 941 1033
rect 959 1028 964 1033
rect 878 1020 883 1025
rect 778 938 783 943
rect 835 939 840 944
rect 669 920 674 925
rect 685 920 690 925
rect 701 920 706 925
rect 717 920 722 925
rect 635 735 640 740
rect 824 735 829 740
rect 982 735 987 740
rect 406 717 411 722
rect 424 717 429 722
rect 690 719 695 724
rect 706 719 711 724
rect 722 719 727 724
rect 738 719 743 724
rect 754 719 759 724
rect 883 719 888 724
rect 899 719 904 724
rect 915 719 920 724
rect 931 719 936 724
rect 212 699 217 704
rect 272 699 277 704
rect 1045 718 1050 723
rect 1061 718 1066 723
rect 1077 718 1082 723
rect 1198 725 1203 730
rect 1221 725 1226 730
rect 1140 717 1145 722
rect 1872 699 1877 704
rect 1895 699 1900 704
rect 323 678 328 683
rect 341 678 346 683
rect 2008 699 2013 704
rect 2031 699 2036 704
rect 2154 701 2159 706
rect 2177 701 2182 706
rect 1953 691 1958 696
rect 2089 691 2094 696
rect 2301 701 2306 706
rect 2324 701 2329 706
rect 2235 693 2240 698
rect 2513 700 2518 705
rect 2536 700 2541 705
rect 2382 693 2387 698
rect 2649 700 2654 705
rect 2672 700 2677 705
rect 2795 702 2800 707
rect 2818 702 2823 707
rect 2594 692 2599 697
rect 2730 692 2735 697
rect 2942 702 2947 707
rect 2965 702 2970 707
rect 2876 694 2881 699
rect 3023 694 3028 699
rect 484 656 489 661
rect 1872 591 1877 596
rect 1895 591 1900 596
rect 2016 591 2021 596
rect 2039 591 2044 596
rect 2165 593 2170 598
rect 2188 593 2193 598
rect 2310 594 2315 599
rect 2333 594 2338 599
rect 1953 583 1958 588
rect 2097 583 2102 588
rect 2246 585 2251 590
rect 2391 586 2396 591
rect 1565 521 1570 526
rect 1588 521 1593 526
rect 403 495 408 500
rect 421 495 426 500
rect 209 477 214 482
rect 269 477 274 482
rect 320 456 325 461
rect 338 456 343 461
rect 751 479 756 484
rect 774 479 779 484
rect 693 471 698 476
rect 898 479 903 484
rect 921 479 926 484
rect 1644 514 1649 519
rect 840 471 845 476
rect 1044 477 1049 482
rect 1067 477 1072 482
rect 986 469 991 474
rect 1180 477 1185 482
rect 1203 477 1208 482
rect 1122 469 1127 474
rect 481 434 486 439
rect 2273 411 2278 416
rect 2296 411 2301 416
rect 742 372 747 377
rect 765 372 770 377
rect 1564 403 1569 408
rect 1587 403 1592 408
rect 684 364 689 369
rect 887 371 892 376
rect 910 371 915 376
rect 1416 375 1421 380
rect 1454 375 1459 380
rect 1643 395 1648 400
rect 829 363 834 368
rect 1036 369 1041 374
rect 1059 369 1064 374
rect 978 361 983 366
rect 1180 369 1185 374
rect 1203 369 1208 374
rect 1122 361 1127 366
rect 2409 411 2414 416
rect 2432 411 2437 416
rect 2555 413 2560 418
rect 2578 413 2583 418
rect 2354 403 2359 408
rect 2490 403 2495 408
rect 2702 413 2707 418
rect 2725 413 2730 418
rect 2636 405 2641 410
rect 2783 405 2788 410
rect 18 304 23 309
rect 2081 342 2086 347
rect 406 310 411 315
rect 424 310 429 315
rect 2012 325 2017 330
rect 2036 325 2041 330
rect 1563 299 1568 304
rect 1586 299 1591 304
rect 2273 303 2278 308
rect 2296 303 2301 308
rect 77 288 82 293
rect 93 288 98 293
rect 109 288 114 293
rect 125 288 130 293
rect 212 292 217 297
rect 272 292 277 297
rect 323 271 328 276
rect 341 271 346 276
rect 1644 291 1649 296
rect 2417 303 2422 308
rect 2440 303 2445 308
rect 2566 305 2571 310
rect 2589 305 2594 310
rect 2711 306 2716 311
rect 2734 306 2739 311
rect 2354 295 2359 300
rect 2498 295 2503 300
rect 2647 297 2652 302
rect 2792 298 2797 303
rect 484 249 489 254
rect 1563 203 1568 208
rect 1586 203 1591 208
rect 1643 195 1648 200
rect 406 135 411 140
rect 424 135 429 140
rect 212 117 217 122
rect 272 117 277 122
rect 323 96 328 101
rect 341 96 346 101
rect 2162 105 2167 110
rect 2180 105 2185 110
rect 2024 87 2029 92
rect 484 74 489 79
rect 2079 66 2084 71
rect 2097 66 2102 71
rect 2240 44 2245 49
rect 1476 -19 1481 -14
rect 1539 -37 1544 -32
rect 1555 -37 1560 -32
rect 1571 -37 1576 -32
rect 2156 -78 2161 -73
rect 2174 -78 2179 -73
rect 2018 -96 2023 -91
rect 1360 -144 1365 -139
rect 1383 -144 1388 -139
rect 2073 -117 2078 -112
rect 2091 -117 2096 -112
rect 1302 -152 1307 -147
rect 1506 -146 1511 -141
rect 1529 -146 1534 -141
rect 1448 -154 1453 -149
rect 1642 -146 1647 -141
rect 1665 -146 1670 -141
rect 1584 -154 1589 -149
rect 2234 -139 2239 -134
rect 1310 -267 1315 -262
rect 1328 -267 1333 -262
rect 2144 -250 2149 -245
rect 2162 -250 2167 -245
rect 1648 -267 1653 -262
rect 1666 -267 1671 -262
rect 2006 -268 2011 -263
rect 1474 -285 1479 -280
rect 1250 -328 1255 -323
rect 1393 -306 1398 -301
rect 1411 -306 1416 -301
rect 1806 -285 1811 -280
rect 2061 -289 2066 -284
rect 2079 -289 2084 -284
rect 1588 -328 1593 -323
rect 1731 -306 1736 -301
rect 1749 -306 1754 -301
rect 2222 -311 2227 -306
rect 2135 -434 2140 -429
rect 2153 -434 2158 -429
rect 1997 -452 2002 -447
rect 2052 -473 2057 -468
rect 2070 -473 2075 -468
rect 2213 -495 2218 -490
<< ptransistor >>
rect 936 1057 941 1062
rect 959 1057 964 1062
rect 878 1042 883 1047
rect 669 956 674 961
rect 685 956 690 961
rect 701 956 706 961
rect 717 956 722 961
rect 778 960 783 965
rect 835 961 840 966
rect 635 757 640 762
rect 690 753 695 758
rect 706 753 711 758
rect 722 753 727 758
rect 738 753 743 758
rect 754 753 759 758
rect 824 757 829 762
rect 212 721 217 726
rect 272 721 277 726
rect 883 753 888 758
rect 899 753 904 758
rect 915 753 920 758
rect 931 753 936 758
rect 982 757 987 762
rect 1045 752 1050 757
rect 1061 752 1066 757
rect 1077 752 1082 757
rect 1198 754 1203 759
rect 1221 754 1226 759
rect 323 717 328 722
rect 341 717 346 722
rect 1140 739 1145 744
rect 1872 728 1877 733
rect 1895 728 1900 733
rect 2008 728 2013 733
rect 2031 728 2036 733
rect 2154 730 2159 735
rect 2177 730 2182 735
rect 2301 730 2306 735
rect 2324 730 2329 735
rect 1953 713 1958 718
rect 2089 713 2094 718
rect 2235 715 2240 720
rect 2513 729 2518 734
rect 2536 729 2541 734
rect 2649 729 2654 734
rect 2672 729 2677 734
rect 2795 731 2800 736
rect 2818 731 2823 736
rect 2942 731 2947 736
rect 2965 731 2970 736
rect 2382 715 2387 720
rect 406 678 411 683
rect 424 678 429 683
rect 484 678 489 683
rect 2594 714 2599 719
rect 2730 714 2735 719
rect 2876 716 2881 721
rect 3023 716 3028 721
rect 1872 620 1877 625
rect 1895 620 1900 625
rect 2016 620 2021 625
rect 2039 620 2044 625
rect 2165 622 2170 627
rect 2188 622 2193 627
rect 2310 623 2315 628
rect 2333 623 2338 628
rect 1953 605 1958 610
rect 2097 605 2102 610
rect 2246 607 2251 612
rect 2391 608 2396 613
rect 1565 550 1570 555
rect 1588 550 1593 555
rect 209 499 214 504
rect 269 499 274 504
rect 1644 536 1649 541
rect 751 508 756 513
rect 774 508 779 513
rect 898 508 903 513
rect 921 508 926 513
rect 320 495 325 500
rect 338 495 343 500
rect 693 493 698 498
rect 840 493 845 498
rect 1044 506 1049 511
rect 1067 506 1072 511
rect 1180 506 1185 511
rect 1203 506 1208 511
rect 986 491 991 496
rect 403 456 408 461
rect 421 456 426 461
rect 481 456 486 461
rect 1122 491 1127 496
rect 2273 440 2278 445
rect 2296 440 2301 445
rect 2409 440 2414 445
rect 2432 440 2437 445
rect 2555 442 2560 447
rect 2578 442 2583 447
rect 2702 442 2707 447
rect 2725 442 2730 447
rect 1564 432 1569 437
rect 1587 432 1592 437
rect 742 401 747 406
rect 765 401 770 406
rect 684 386 689 391
rect 887 400 892 405
rect 910 400 915 405
rect 1643 417 1648 422
rect 2354 425 2359 430
rect 2490 425 2495 430
rect 2636 427 2641 432
rect 2783 427 2788 432
rect 829 385 834 390
rect 1036 398 1041 403
rect 1059 398 1064 403
rect 1180 398 1185 403
rect 1203 398 1208 403
rect 978 383 983 388
rect 1122 383 1127 388
rect 1416 397 1421 402
rect 1454 397 1459 402
rect 18 326 23 331
rect 2012 362 2017 367
rect 2036 362 2041 367
rect 2081 364 2086 369
rect 77 322 82 327
rect 93 322 98 327
rect 109 322 114 327
rect 125 322 130 327
rect 212 314 217 319
rect 272 314 277 319
rect 1563 328 1568 333
rect 1586 328 1591 333
rect 2273 332 2278 337
rect 2296 332 2301 337
rect 2417 332 2422 337
rect 2440 332 2445 337
rect 2566 334 2571 339
rect 2589 334 2594 339
rect 2711 335 2716 340
rect 2734 335 2739 340
rect 323 310 328 315
rect 341 310 346 315
rect 1644 313 1649 318
rect 2354 317 2359 322
rect 2498 317 2503 322
rect 2647 319 2652 324
rect 2792 320 2797 325
rect 406 271 411 276
rect 424 271 429 276
rect 484 271 489 276
rect 1563 232 1568 237
rect 1586 232 1591 237
rect 1643 217 1648 222
rect 212 139 217 144
rect 272 139 277 144
rect 323 135 328 140
rect 341 135 346 140
rect 2024 109 2029 114
rect 406 96 411 101
rect 424 96 429 101
rect 484 96 489 101
rect 2079 105 2084 110
rect 2097 105 2102 110
rect 2162 66 2167 71
rect 2180 66 2185 71
rect 2240 66 2245 71
rect 1476 3 1481 8
rect 1539 -1 1544 4
rect 1555 -1 1560 4
rect 1571 -1 1576 4
rect 2018 -74 2023 -69
rect 2073 -78 2078 -73
rect 2091 -78 2096 -73
rect 1360 -115 1365 -110
rect 1383 -115 1388 -110
rect 1302 -130 1307 -125
rect 1506 -117 1511 -112
rect 1529 -117 1534 -112
rect 1642 -117 1647 -112
rect 1665 -117 1670 -112
rect 1448 -132 1453 -127
rect 1584 -132 1589 -127
rect 2156 -117 2161 -112
rect 2174 -117 2179 -112
rect 2234 -117 2239 -112
rect 1393 -267 1398 -262
rect 1411 -267 1416 -262
rect 1474 -263 1479 -258
rect 2006 -246 2011 -241
rect 2061 -250 2066 -245
rect 2079 -250 2084 -245
rect 1731 -267 1736 -262
rect 1749 -267 1754 -262
rect 1806 -263 1811 -258
rect 1250 -306 1255 -301
rect 1310 -306 1315 -301
rect 1328 -306 1333 -301
rect 1588 -306 1593 -301
rect 1648 -306 1653 -301
rect 1666 -306 1671 -301
rect 2144 -289 2149 -284
rect 2162 -289 2167 -284
rect 2222 -289 2227 -284
rect 1997 -430 2002 -425
rect 2052 -434 2057 -429
rect 2070 -434 2075 -429
rect 2135 -473 2140 -468
rect 2153 -473 2158 -468
rect 2213 -473 2218 -468
<< ndiffusion >>
rect 934 1028 936 1033
rect 941 1028 943 1033
rect 957 1028 959 1033
rect 964 1028 966 1033
rect 875 1020 878 1025
rect 883 1020 885 1025
rect 776 938 778 943
rect 783 938 786 943
rect 833 939 835 944
rect 840 939 843 944
rect 666 920 669 925
rect 674 920 677 925
rect 682 920 685 925
rect 690 920 693 925
rect 698 920 701 925
rect 706 920 709 925
rect 714 920 717 925
rect 722 920 725 925
rect 632 735 635 740
rect 640 735 642 740
rect 821 735 824 740
rect 829 735 831 740
rect 979 735 982 740
rect 987 735 989 740
rect 403 717 406 722
rect 411 717 424 722
rect 429 717 432 722
rect 687 719 690 724
rect 695 719 706 724
rect 711 719 722 724
rect 727 719 738 724
rect 743 719 754 724
rect 759 719 762 724
rect 881 719 883 724
rect 888 719 899 724
rect 904 719 915 724
rect 920 719 931 724
rect 936 719 939 724
rect 210 699 212 704
rect 217 699 220 704
rect 269 699 272 704
rect 277 699 279 704
rect 1039 718 1045 723
rect 1050 718 1061 723
rect 1066 718 1077 723
rect 1082 718 1085 723
rect 1196 725 1198 730
rect 1203 725 1205 730
rect 1219 725 1221 730
rect 1226 725 1228 730
rect 1137 717 1140 722
rect 1145 717 1147 722
rect 1870 699 1872 704
rect 1877 699 1879 704
rect 1893 699 1895 704
rect 1900 699 1902 704
rect 320 678 323 683
rect 328 678 341 683
rect 346 678 349 683
rect 2006 699 2008 704
rect 2013 699 2015 704
rect 2029 699 2031 704
rect 2036 699 2038 704
rect 2152 701 2154 706
rect 2159 701 2161 706
rect 2175 701 2177 706
rect 2182 701 2184 706
rect 1951 691 1953 696
rect 1958 691 1961 696
rect 2087 691 2089 696
rect 2094 691 2097 696
rect 2299 701 2301 706
rect 2306 701 2308 706
rect 2322 701 2324 706
rect 2329 701 2331 706
rect 2233 693 2235 698
rect 2240 693 2243 698
rect 2511 700 2513 705
rect 2518 700 2520 705
rect 2534 700 2536 705
rect 2541 700 2543 705
rect 2380 693 2382 698
rect 2387 693 2390 698
rect 2647 700 2649 705
rect 2654 700 2656 705
rect 2670 700 2672 705
rect 2677 700 2679 705
rect 2793 702 2795 707
rect 2800 702 2802 707
rect 2816 702 2818 707
rect 2823 702 2825 707
rect 2592 692 2594 697
rect 2599 692 2602 697
rect 2728 692 2730 697
rect 2735 692 2738 697
rect 2940 702 2942 707
rect 2947 702 2949 707
rect 2963 702 2965 707
rect 2970 702 2972 707
rect 2874 694 2876 699
rect 2881 694 2884 699
rect 3021 694 3023 699
rect 3028 694 3031 699
rect 482 656 484 661
rect 489 656 492 661
rect 1870 591 1872 596
rect 1877 591 1879 596
rect 1893 591 1895 596
rect 1900 591 1902 596
rect 2014 591 2016 596
rect 2021 591 2023 596
rect 2037 591 2039 596
rect 2044 591 2046 596
rect 2163 593 2165 598
rect 2170 593 2172 598
rect 2186 593 2188 598
rect 2193 593 2195 598
rect 2308 594 2310 599
rect 2315 594 2317 599
rect 2331 594 2333 599
rect 2338 594 2340 599
rect 1951 583 1953 588
rect 1958 583 1961 588
rect 2095 583 2097 588
rect 2102 583 2105 588
rect 2244 585 2246 590
rect 2251 585 2254 590
rect 2389 586 2391 591
rect 2396 586 2399 591
rect 1563 521 1565 526
rect 1570 521 1572 526
rect 1586 521 1588 526
rect 1593 521 1595 526
rect 400 495 403 500
rect 408 495 421 500
rect 426 495 429 500
rect 207 477 209 482
rect 214 477 217 482
rect 266 477 269 482
rect 274 477 276 482
rect 317 456 320 461
rect 325 456 338 461
rect 343 456 346 461
rect 749 479 751 484
rect 756 479 758 484
rect 772 479 774 484
rect 779 479 781 484
rect 690 471 693 476
rect 698 471 700 476
rect 896 479 898 484
rect 903 479 905 484
rect 919 479 921 484
rect 926 479 928 484
rect 1642 514 1644 519
rect 1649 514 1652 519
rect 837 471 840 476
rect 845 471 847 476
rect 1042 477 1044 482
rect 1049 477 1051 482
rect 1065 477 1067 482
rect 1072 477 1074 482
rect 983 469 986 474
rect 991 469 993 474
rect 1178 477 1180 482
rect 1185 477 1187 482
rect 1201 477 1203 482
rect 1208 477 1210 482
rect 1119 469 1122 474
rect 1127 469 1129 474
rect 479 434 481 439
rect 486 434 489 439
rect 2271 411 2273 416
rect 2278 411 2280 416
rect 2294 411 2296 416
rect 2301 411 2303 416
rect 740 372 742 377
rect 747 372 749 377
rect 763 372 765 377
rect 770 372 772 377
rect 1562 403 1564 408
rect 1569 403 1571 408
rect 1585 403 1587 408
rect 1592 403 1594 408
rect 681 364 684 369
rect 689 364 691 369
rect 885 371 887 376
rect 892 371 894 376
rect 908 371 910 376
rect 915 371 917 376
rect 1414 375 1416 380
rect 1421 375 1424 380
rect 1452 375 1454 380
rect 1459 375 1462 380
rect 1641 395 1643 400
rect 1648 395 1651 400
rect 826 363 829 368
rect 834 363 836 368
rect 1034 369 1036 374
rect 1041 369 1043 374
rect 1057 369 1059 374
rect 1064 369 1066 374
rect 975 361 978 366
rect 983 361 985 366
rect 1178 369 1180 374
rect 1185 369 1187 374
rect 1201 369 1203 374
rect 1208 369 1210 374
rect 1119 361 1122 366
rect 1127 361 1129 366
rect 2407 411 2409 416
rect 2414 411 2416 416
rect 2430 411 2432 416
rect 2437 411 2439 416
rect 2553 413 2555 418
rect 2560 413 2562 418
rect 2576 413 2578 418
rect 2583 413 2585 418
rect 2352 403 2354 408
rect 2359 403 2362 408
rect 2488 403 2490 408
rect 2495 403 2498 408
rect 2700 413 2702 418
rect 2707 413 2709 418
rect 2723 413 2725 418
rect 2730 413 2732 418
rect 2634 405 2636 410
rect 2641 405 2644 410
rect 2781 405 2783 410
rect 2788 405 2791 410
rect 15 304 18 309
rect 23 304 25 309
rect 2079 342 2081 347
rect 2086 342 2089 347
rect 403 310 406 315
rect 411 310 424 315
rect 429 310 432 315
rect 2010 325 2012 330
rect 2017 325 2023 330
rect 2028 325 2036 330
rect 2041 325 2043 330
rect 1561 299 1563 304
rect 1568 299 1570 304
rect 1584 299 1586 304
rect 1591 299 1593 304
rect 2271 303 2273 308
rect 2278 303 2280 308
rect 2294 303 2296 308
rect 2301 303 2303 308
rect 75 288 77 293
rect 82 288 93 293
rect 98 288 109 293
rect 114 288 125 293
rect 130 288 133 293
rect 210 292 212 297
rect 217 292 220 297
rect 269 292 272 297
rect 277 292 279 297
rect 320 271 323 276
rect 328 271 341 276
rect 346 271 349 276
rect 1642 291 1644 296
rect 1649 291 1652 296
rect 2415 303 2417 308
rect 2422 303 2424 308
rect 2438 303 2440 308
rect 2445 303 2447 308
rect 2564 305 2566 310
rect 2571 305 2573 310
rect 2587 305 2589 310
rect 2594 305 2596 310
rect 2709 306 2711 311
rect 2716 306 2718 311
rect 2732 306 2734 311
rect 2739 306 2741 311
rect 2352 295 2354 300
rect 2359 295 2362 300
rect 2496 295 2498 300
rect 2503 295 2506 300
rect 2645 297 2647 302
rect 2652 297 2655 302
rect 2790 298 2792 303
rect 2797 298 2800 303
rect 482 249 484 254
rect 489 249 492 254
rect 1561 203 1563 208
rect 1568 203 1570 208
rect 1584 203 1586 208
rect 1591 203 1593 208
rect 1641 195 1643 200
rect 1648 195 1651 200
rect 403 135 406 140
rect 411 135 424 140
rect 429 135 432 140
rect 210 117 212 122
rect 217 117 220 122
rect 269 117 272 122
rect 277 117 279 122
rect 320 96 323 101
rect 328 96 341 101
rect 346 96 349 101
rect 2159 105 2162 110
rect 2167 105 2180 110
rect 2185 105 2188 110
rect 2021 87 2024 92
rect 2029 87 2031 92
rect 482 74 484 79
rect 489 74 492 79
rect 2076 66 2079 71
rect 2084 66 2097 71
rect 2102 66 2105 71
rect 2238 44 2240 49
rect 2245 44 2248 49
rect 1473 -19 1476 -14
rect 1481 -19 1483 -14
rect 1536 -37 1539 -32
rect 1544 -37 1547 -32
rect 1552 -37 1555 -32
rect 1560 -37 1563 -32
rect 1568 -37 1571 -32
rect 1576 -37 1579 -32
rect 2153 -78 2156 -73
rect 2161 -78 2174 -73
rect 2179 -78 2182 -73
rect 2015 -96 2018 -91
rect 2023 -96 2025 -91
rect 1358 -144 1360 -139
rect 1365 -144 1367 -139
rect 1381 -144 1383 -139
rect 1388 -144 1390 -139
rect 2070 -117 2073 -112
rect 2078 -117 2091 -112
rect 2096 -117 2099 -112
rect 1299 -152 1302 -147
rect 1307 -152 1309 -147
rect 1504 -146 1506 -141
rect 1511 -146 1513 -141
rect 1527 -146 1529 -141
rect 1534 -146 1536 -141
rect 1445 -154 1448 -149
rect 1453 -154 1455 -149
rect 1640 -146 1642 -141
rect 1647 -146 1649 -141
rect 1663 -146 1665 -141
rect 1670 -146 1672 -141
rect 1581 -154 1584 -149
rect 1589 -154 1591 -149
rect 2232 -139 2234 -134
rect 2239 -139 2242 -134
rect 1307 -267 1310 -262
rect 1315 -267 1328 -262
rect 1333 -267 1336 -262
rect 2141 -250 2144 -245
rect 2149 -250 2162 -245
rect 2167 -250 2170 -245
rect 1645 -267 1648 -262
rect 1653 -267 1666 -262
rect 1671 -267 1674 -262
rect 2003 -268 2006 -263
rect 2011 -268 2013 -263
rect 1472 -285 1474 -280
rect 1479 -285 1482 -280
rect 1247 -328 1250 -323
rect 1255 -328 1257 -323
rect 1390 -306 1393 -301
rect 1398 -306 1411 -301
rect 1416 -306 1419 -301
rect 1804 -285 1806 -280
rect 1811 -285 1814 -280
rect 2058 -289 2061 -284
rect 2066 -289 2079 -284
rect 2084 -289 2087 -284
rect 1585 -328 1588 -323
rect 1593 -328 1595 -323
rect 1728 -306 1731 -301
rect 1736 -306 1749 -301
rect 1754 -306 1757 -301
rect 2220 -311 2222 -306
rect 2227 -311 2230 -306
rect 2132 -434 2135 -429
rect 2140 -434 2153 -429
rect 2158 -434 2161 -429
rect 1994 -452 1997 -447
rect 2002 -452 2004 -447
rect 2049 -473 2052 -468
rect 2057 -473 2070 -468
rect 2075 -473 2078 -468
rect 2211 -495 2213 -490
rect 2218 -495 2221 -490
<< pdiffusion >>
rect 934 1057 936 1062
rect 941 1057 947 1062
rect 952 1057 959 1062
rect 964 1057 966 1062
rect 875 1042 878 1047
rect 883 1042 885 1047
rect 666 956 669 961
rect 674 956 685 961
rect 690 956 701 961
rect 706 956 717 961
rect 722 956 725 961
rect 776 960 778 965
rect 783 960 786 965
rect 833 961 835 966
rect 840 961 843 966
rect 632 757 635 762
rect 640 757 642 762
rect 687 753 690 758
rect 695 753 698 758
rect 703 753 706 758
rect 711 753 714 758
rect 719 753 722 758
rect 727 753 730 758
rect 735 753 738 758
rect 743 753 746 758
rect 751 753 754 758
rect 759 753 762 758
rect 821 757 824 762
rect 829 757 831 762
rect 210 721 212 726
rect 217 721 220 726
rect 269 721 272 726
rect 277 721 279 726
rect 880 753 883 758
rect 888 753 891 758
rect 896 753 899 758
rect 904 753 907 758
rect 912 753 915 758
rect 920 753 923 758
rect 928 753 931 758
rect 936 753 939 758
rect 979 757 982 762
rect 987 757 989 762
rect 1042 752 1045 757
rect 1050 752 1053 757
rect 1058 752 1061 757
rect 1066 752 1069 757
rect 1074 752 1077 757
rect 1082 752 1085 757
rect 1196 754 1198 759
rect 1203 754 1209 759
rect 1214 754 1221 759
rect 1226 754 1228 759
rect 320 717 323 722
rect 328 717 341 722
rect 346 717 349 722
rect 1137 739 1140 744
rect 1145 739 1147 744
rect 1870 728 1872 733
rect 1877 728 1884 733
rect 1889 728 1895 733
rect 1900 728 1902 733
rect 2006 728 2008 733
rect 2013 728 2020 733
rect 2025 728 2031 733
rect 2036 728 2038 733
rect 2152 730 2154 735
rect 2159 730 2166 735
rect 2171 730 2177 735
rect 2182 730 2184 735
rect 2299 730 2301 735
rect 2306 730 2313 735
rect 2318 730 2324 735
rect 2329 730 2331 735
rect 1951 713 1953 718
rect 1958 713 1961 718
rect 2087 713 2089 718
rect 2094 713 2097 718
rect 2233 715 2235 720
rect 2240 715 2243 720
rect 2511 729 2513 734
rect 2518 729 2525 734
rect 2530 729 2536 734
rect 2541 729 2543 734
rect 2647 729 2649 734
rect 2654 729 2661 734
rect 2666 729 2672 734
rect 2677 729 2679 734
rect 2793 731 2795 736
rect 2800 731 2807 736
rect 2812 731 2818 736
rect 2823 731 2825 736
rect 2940 731 2942 736
rect 2947 731 2954 736
rect 2959 731 2965 736
rect 2970 731 2972 736
rect 2380 715 2382 720
rect 2387 715 2390 720
rect 403 678 406 683
rect 411 678 424 683
rect 429 678 432 683
rect 482 678 484 683
rect 489 678 492 683
rect 2592 714 2594 719
rect 2599 714 2602 719
rect 2728 714 2730 719
rect 2735 714 2738 719
rect 2874 716 2876 721
rect 2881 716 2884 721
rect 3021 716 3023 721
rect 3028 716 3031 721
rect 1870 620 1872 625
rect 1877 620 1884 625
rect 1889 620 1895 625
rect 1900 620 1902 625
rect 2014 620 2016 625
rect 2021 620 2028 625
rect 2033 620 2039 625
rect 2044 620 2046 625
rect 2163 622 2165 627
rect 2170 622 2177 627
rect 2182 622 2188 627
rect 2193 622 2195 627
rect 2308 623 2310 628
rect 2315 623 2322 628
rect 2327 623 2333 628
rect 2338 623 2340 628
rect 1951 605 1953 610
rect 1958 605 1961 610
rect 2095 605 2097 610
rect 2102 605 2105 610
rect 2244 607 2246 612
rect 2251 607 2254 612
rect 2389 608 2391 613
rect 2396 608 2399 613
rect 1563 550 1565 555
rect 1570 550 1577 555
rect 1582 550 1588 555
rect 1593 550 1595 555
rect 207 499 209 504
rect 214 499 217 504
rect 266 499 269 504
rect 274 499 276 504
rect 1642 536 1644 541
rect 1649 536 1652 541
rect 749 508 751 513
rect 756 508 762 513
rect 767 508 774 513
rect 779 508 781 513
rect 896 508 898 513
rect 903 508 909 513
rect 914 508 921 513
rect 926 508 928 513
rect 317 495 320 500
rect 325 495 338 500
rect 343 495 346 500
rect 690 493 693 498
rect 698 493 700 498
rect 837 493 840 498
rect 845 493 847 498
rect 1042 506 1044 511
rect 1049 506 1055 511
rect 1060 506 1067 511
rect 1072 506 1074 511
rect 1178 506 1180 511
rect 1185 506 1191 511
rect 1196 506 1203 511
rect 1208 506 1210 511
rect 983 491 986 496
rect 991 491 993 496
rect 400 456 403 461
rect 408 456 421 461
rect 426 456 429 461
rect 479 456 481 461
rect 486 456 489 461
rect 1119 491 1122 496
rect 1127 491 1129 496
rect 2271 440 2273 445
rect 2278 440 2285 445
rect 2290 440 2296 445
rect 2301 440 2303 445
rect 2407 440 2409 445
rect 2414 440 2421 445
rect 2426 440 2432 445
rect 2437 440 2439 445
rect 2553 442 2555 447
rect 2560 442 2567 447
rect 2572 442 2578 447
rect 2583 442 2585 447
rect 2700 442 2702 447
rect 2707 442 2714 447
rect 2719 442 2725 447
rect 2730 442 2732 447
rect 1562 432 1564 437
rect 1569 432 1576 437
rect 1581 432 1587 437
rect 1592 432 1594 437
rect 740 401 742 406
rect 747 401 753 406
rect 758 401 765 406
rect 770 401 772 406
rect 681 386 684 391
rect 689 386 691 391
rect 885 400 887 405
rect 892 400 898 405
rect 903 400 910 405
rect 915 400 917 405
rect 1641 417 1643 422
rect 1648 417 1651 422
rect 2352 425 2354 430
rect 2359 425 2362 430
rect 2488 425 2490 430
rect 2495 425 2498 430
rect 2634 427 2636 432
rect 2641 427 2644 432
rect 2781 427 2783 432
rect 2788 427 2791 432
rect 826 385 829 390
rect 834 385 836 390
rect 1034 398 1036 403
rect 1041 398 1047 403
rect 1052 398 1059 403
rect 1064 398 1066 403
rect 1178 398 1180 403
rect 1185 398 1191 403
rect 1196 398 1203 403
rect 1208 398 1210 403
rect 975 383 978 388
rect 983 383 985 388
rect 1119 383 1122 388
rect 1127 383 1129 388
rect 1414 397 1416 402
rect 1421 397 1424 402
rect 1452 397 1454 402
rect 1459 397 1462 402
rect 15 326 18 331
rect 23 326 25 331
rect 2010 362 2012 367
rect 2017 362 2019 367
rect 2034 362 2036 367
rect 2041 362 2043 367
rect 2079 364 2081 369
rect 2086 364 2089 369
rect 74 322 77 327
rect 82 322 85 327
rect 90 322 93 327
rect 98 322 101 327
rect 106 322 109 327
rect 114 322 117 327
rect 122 322 125 327
rect 130 322 133 327
rect 210 314 212 319
rect 217 314 220 319
rect 269 314 272 319
rect 277 314 279 319
rect 1561 328 1563 333
rect 1568 328 1575 333
rect 1580 328 1586 333
rect 1591 328 1593 333
rect 2271 332 2273 337
rect 2278 332 2285 337
rect 2290 332 2296 337
rect 2301 332 2303 337
rect 2415 332 2417 337
rect 2422 332 2429 337
rect 2434 332 2440 337
rect 2445 332 2447 337
rect 2564 334 2566 339
rect 2571 334 2578 339
rect 2583 334 2589 339
rect 2594 334 2596 339
rect 2709 335 2711 340
rect 2716 335 2723 340
rect 2728 335 2734 340
rect 2739 335 2741 340
rect 320 310 323 315
rect 328 310 341 315
rect 346 310 349 315
rect 1642 313 1644 318
rect 1649 313 1652 318
rect 2352 317 2354 322
rect 2359 317 2362 322
rect 2496 317 2498 322
rect 2503 317 2506 322
rect 2645 319 2647 324
rect 2652 319 2655 324
rect 2790 320 2792 325
rect 2797 320 2800 325
rect 403 271 406 276
rect 411 271 424 276
rect 429 271 432 276
rect 482 271 484 276
rect 489 271 492 276
rect 1561 232 1563 237
rect 1568 232 1575 237
rect 1580 232 1586 237
rect 1591 232 1593 237
rect 1641 217 1643 222
rect 1648 217 1651 222
rect 210 139 212 144
rect 217 139 220 144
rect 269 139 272 144
rect 277 139 279 144
rect 320 135 323 140
rect 328 135 341 140
rect 346 135 349 140
rect 2021 109 2024 114
rect 2029 109 2031 114
rect 403 96 406 101
rect 411 96 424 101
rect 429 96 432 101
rect 482 96 484 101
rect 489 96 492 101
rect 2076 105 2079 110
rect 2084 105 2097 110
rect 2102 105 2105 110
rect 2159 66 2162 71
rect 2167 66 2180 71
rect 2185 66 2188 71
rect 2238 66 2240 71
rect 2245 66 2248 71
rect 1473 3 1476 8
rect 1481 3 1483 8
rect 1536 -1 1539 4
rect 1544 -1 1555 4
rect 1560 -1 1571 4
rect 1576 -1 1579 4
rect 2015 -74 2018 -69
rect 2023 -74 2025 -69
rect 2070 -78 2073 -73
rect 2078 -78 2091 -73
rect 2096 -78 2099 -73
rect 1358 -115 1360 -110
rect 1365 -115 1371 -110
rect 1376 -115 1383 -110
rect 1388 -115 1390 -110
rect 1299 -130 1302 -125
rect 1307 -130 1309 -125
rect 1504 -117 1506 -112
rect 1511 -117 1517 -112
rect 1522 -117 1529 -112
rect 1534 -117 1536 -112
rect 1640 -117 1642 -112
rect 1647 -117 1653 -112
rect 1658 -117 1665 -112
rect 1670 -117 1672 -112
rect 1445 -132 1448 -127
rect 1453 -132 1455 -127
rect 1581 -132 1584 -127
rect 1589 -132 1591 -127
rect 2153 -117 2156 -112
rect 2161 -117 2174 -112
rect 2179 -117 2182 -112
rect 2232 -117 2234 -112
rect 2239 -117 2242 -112
rect 1390 -267 1393 -262
rect 1398 -267 1411 -262
rect 1416 -267 1419 -262
rect 1472 -263 1474 -258
rect 1479 -263 1482 -258
rect 2003 -246 2006 -241
rect 2011 -246 2013 -241
rect 2058 -250 2061 -245
rect 2066 -250 2079 -245
rect 2084 -250 2087 -245
rect 1728 -267 1731 -262
rect 1736 -267 1749 -262
rect 1754 -267 1757 -262
rect 1804 -263 1806 -258
rect 1811 -263 1814 -258
rect 1247 -306 1250 -301
rect 1255 -306 1257 -301
rect 1307 -306 1310 -301
rect 1315 -306 1328 -301
rect 1333 -306 1336 -301
rect 1585 -306 1588 -301
rect 1593 -306 1595 -301
rect 1645 -306 1648 -301
rect 1653 -306 1666 -301
rect 1671 -306 1674 -301
rect 2141 -289 2144 -284
rect 2149 -289 2162 -284
rect 2167 -289 2170 -284
rect 2220 -289 2222 -284
rect 2227 -289 2230 -284
rect 1994 -430 1997 -425
rect 2002 -430 2004 -425
rect 2049 -434 2052 -429
rect 2057 -434 2070 -429
rect 2075 -434 2078 -429
rect 2132 -473 2135 -468
rect 2140 -473 2153 -468
rect 2158 -473 2161 -468
rect 2211 -473 2213 -468
rect 2218 -473 2221 -468
<< ndcontact >>
rect 929 1028 934 1033
rect 943 1028 947 1033
rect 953 1028 957 1033
rect 966 1028 971 1033
rect 870 1020 875 1025
rect 885 1020 890 1025
rect 771 938 776 943
rect 786 938 791 943
rect 828 939 833 944
rect 843 939 848 944
rect 661 920 666 925
rect 677 920 682 925
rect 693 920 698 925
rect 709 920 714 925
rect 725 920 730 925
rect 627 735 632 740
rect 642 735 647 740
rect 816 735 821 740
rect 831 735 836 740
rect 974 735 979 740
rect 989 735 994 740
rect 398 717 403 722
rect 432 717 437 722
rect 682 719 687 724
rect 762 719 767 724
rect 876 719 881 724
rect 939 719 944 724
rect 205 699 210 704
rect 220 699 225 704
rect 264 699 269 704
rect 279 699 284 704
rect 1034 718 1039 723
rect 1085 718 1090 723
rect 1191 725 1196 730
rect 1205 725 1209 730
rect 1215 725 1219 730
rect 1228 725 1233 730
rect 1132 717 1137 722
rect 1147 717 1152 722
rect 1865 699 1870 704
rect 1879 699 1883 704
rect 1889 699 1893 704
rect 1902 699 1907 704
rect 315 678 320 683
rect 349 678 354 683
rect 2001 699 2006 704
rect 2015 699 2019 704
rect 2025 699 2029 704
rect 2038 699 2043 704
rect 2147 701 2152 706
rect 2161 701 2165 706
rect 2171 701 2175 706
rect 2184 701 2189 706
rect 1946 691 1951 696
rect 1961 691 1966 696
rect 2082 691 2087 696
rect 2097 691 2102 696
rect 2294 701 2299 706
rect 2308 701 2312 706
rect 2318 701 2322 706
rect 2331 701 2336 706
rect 2228 693 2233 698
rect 2243 693 2248 698
rect 2506 700 2511 705
rect 2520 700 2524 705
rect 2530 700 2534 705
rect 2543 700 2548 705
rect 2375 693 2380 698
rect 2390 693 2395 698
rect 2642 700 2647 705
rect 2656 700 2660 705
rect 2666 700 2670 705
rect 2679 700 2684 705
rect 2788 702 2793 707
rect 2802 702 2806 707
rect 2812 702 2816 707
rect 2825 702 2830 707
rect 2587 692 2592 697
rect 2602 692 2607 697
rect 2723 692 2728 697
rect 2738 692 2743 697
rect 2935 702 2940 707
rect 2949 702 2953 707
rect 2959 702 2963 707
rect 2972 702 2977 707
rect 2869 694 2874 699
rect 2884 694 2889 699
rect 3016 694 3021 699
rect 3031 694 3036 699
rect 477 656 482 661
rect 492 656 497 661
rect 1865 591 1870 596
rect 1879 591 1883 596
rect 1889 591 1893 596
rect 1902 591 1907 596
rect 2009 591 2014 596
rect 2023 591 2027 596
rect 2033 591 2037 596
rect 2046 591 2051 596
rect 2158 593 2163 598
rect 2172 593 2176 598
rect 2182 593 2186 598
rect 2195 593 2200 598
rect 2303 594 2308 599
rect 2317 594 2321 599
rect 2327 594 2331 599
rect 2340 594 2345 599
rect 1946 583 1951 588
rect 1961 583 1966 588
rect 2090 583 2095 588
rect 2105 583 2110 588
rect 2239 585 2244 590
rect 2254 585 2259 590
rect 2384 586 2389 591
rect 2399 586 2404 591
rect 1558 521 1563 526
rect 1572 521 1576 526
rect 1582 521 1586 526
rect 1595 521 1600 526
rect 395 495 400 500
rect 429 495 434 500
rect 202 477 207 482
rect 217 477 222 482
rect 261 477 266 482
rect 276 477 281 482
rect 312 456 317 461
rect 346 456 351 461
rect 744 479 749 484
rect 758 479 762 484
rect 768 479 772 484
rect 781 479 786 484
rect 685 471 690 476
rect 700 471 705 476
rect 891 479 896 484
rect 905 479 909 484
rect 915 479 919 484
rect 928 479 933 484
rect 1637 514 1642 519
rect 1652 514 1657 519
rect 832 471 837 476
rect 847 471 852 476
rect 1037 477 1042 482
rect 1051 477 1055 482
rect 1061 477 1065 482
rect 1074 477 1079 482
rect 978 469 983 474
rect 993 469 998 474
rect 1173 477 1178 482
rect 1187 477 1191 482
rect 1197 477 1201 482
rect 1210 477 1215 482
rect 1114 469 1119 474
rect 1129 469 1134 474
rect 474 434 479 439
rect 489 434 494 439
rect 2266 411 2271 416
rect 2280 411 2284 416
rect 2290 411 2294 416
rect 2303 411 2308 416
rect 735 372 740 377
rect 749 372 753 377
rect 759 372 763 377
rect 772 372 777 377
rect 1557 403 1562 408
rect 1571 403 1575 408
rect 1581 403 1585 408
rect 1594 403 1599 408
rect 676 364 681 369
rect 691 364 696 369
rect 880 371 885 376
rect 894 371 898 376
rect 904 371 908 376
rect 917 371 922 376
rect 1409 375 1414 380
rect 1424 375 1429 380
rect 1447 375 1452 380
rect 1462 375 1467 380
rect 1636 395 1641 400
rect 1651 395 1656 400
rect 821 363 826 368
rect 836 363 841 368
rect 1029 369 1034 374
rect 1043 369 1047 374
rect 1053 369 1057 374
rect 1066 369 1071 374
rect 970 361 975 366
rect 985 361 990 366
rect 1173 369 1178 374
rect 1187 369 1191 374
rect 1197 369 1201 374
rect 1210 369 1215 374
rect 1114 361 1119 366
rect 1129 361 1134 366
rect 2402 411 2407 416
rect 2416 411 2420 416
rect 2426 411 2430 416
rect 2439 411 2444 416
rect 2548 413 2553 418
rect 2562 413 2566 418
rect 2572 413 2576 418
rect 2585 413 2590 418
rect 2347 403 2352 408
rect 2362 403 2367 408
rect 2483 403 2488 408
rect 2498 403 2503 408
rect 2695 413 2700 418
rect 2709 413 2713 418
rect 2719 413 2723 418
rect 2732 413 2737 418
rect 2629 405 2634 410
rect 2644 405 2649 410
rect 2776 405 2781 410
rect 2791 405 2796 410
rect 10 304 15 309
rect 25 304 30 309
rect 2074 342 2079 347
rect 2089 342 2094 347
rect 398 310 403 315
rect 432 310 437 315
rect 2005 325 2010 330
rect 2023 325 2028 330
rect 2043 325 2048 330
rect 1556 299 1561 304
rect 1570 299 1574 304
rect 1580 299 1584 304
rect 1593 299 1598 304
rect 2266 303 2271 308
rect 2280 303 2284 308
rect 2290 303 2294 308
rect 2303 303 2308 308
rect 70 288 75 293
rect 133 288 138 293
rect 205 292 210 297
rect 220 292 225 297
rect 264 292 269 297
rect 279 292 284 297
rect 315 271 320 276
rect 349 271 354 276
rect 1637 291 1642 296
rect 1652 291 1657 296
rect 2410 303 2415 308
rect 2424 303 2428 308
rect 2434 303 2438 308
rect 2447 303 2452 308
rect 2559 305 2564 310
rect 2573 305 2577 310
rect 2583 305 2587 310
rect 2596 305 2601 310
rect 2704 306 2709 311
rect 2718 306 2722 311
rect 2728 306 2732 311
rect 2741 306 2746 311
rect 2347 295 2352 300
rect 2362 295 2367 300
rect 2491 295 2496 300
rect 2506 295 2511 300
rect 2640 297 2645 302
rect 2655 297 2660 302
rect 2785 298 2790 303
rect 2800 298 2805 303
rect 477 249 482 254
rect 492 249 497 254
rect 1556 203 1561 208
rect 1570 203 1574 208
rect 1580 203 1584 208
rect 1593 203 1598 208
rect 1636 195 1641 200
rect 1651 195 1656 200
rect 398 135 403 140
rect 432 135 437 140
rect 205 117 210 122
rect 220 117 225 122
rect 264 117 269 122
rect 279 117 284 122
rect 315 96 320 101
rect 349 96 354 101
rect 2154 105 2159 110
rect 2188 105 2193 110
rect 2016 87 2021 92
rect 2031 87 2036 92
rect 477 74 482 79
rect 492 74 497 79
rect 2071 66 2076 71
rect 2105 66 2110 71
rect 2233 44 2238 49
rect 2248 44 2253 49
rect 1468 -19 1473 -14
rect 1483 -19 1488 -14
rect 1531 -37 1536 -32
rect 1547 -37 1552 -32
rect 1563 -37 1568 -32
rect 1579 -37 1584 -32
rect 2148 -78 2153 -73
rect 2182 -78 2187 -73
rect 2010 -96 2015 -91
rect 2025 -96 2030 -91
rect 1353 -144 1358 -139
rect 1367 -144 1371 -139
rect 1377 -144 1381 -139
rect 1390 -144 1395 -139
rect 2065 -117 2070 -112
rect 2099 -117 2104 -112
rect 1294 -152 1299 -147
rect 1309 -152 1314 -147
rect 1499 -146 1504 -141
rect 1513 -146 1517 -141
rect 1523 -146 1527 -141
rect 1536 -146 1541 -141
rect 1440 -154 1445 -149
rect 1455 -154 1460 -149
rect 1635 -146 1640 -141
rect 1649 -146 1653 -141
rect 1659 -146 1663 -141
rect 1672 -146 1677 -141
rect 1576 -154 1581 -149
rect 1591 -154 1596 -149
rect 2227 -139 2232 -134
rect 2242 -139 2247 -134
rect 1302 -267 1307 -262
rect 1336 -267 1341 -262
rect 2136 -250 2141 -245
rect 2170 -250 2175 -245
rect 1640 -267 1645 -262
rect 1674 -267 1679 -262
rect 1998 -268 2003 -263
rect 2013 -268 2018 -263
rect 1467 -285 1472 -280
rect 1482 -285 1487 -280
rect 1242 -328 1247 -323
rect 1257 -328 1262 -323
rect 1385 -306 1390 -301
rect 1419 -306 1424 -301
rect 1799 -285 1804 -280
rect 1814 -285 1819 -280
rect 2053 -289 2058 -284
rect 2087 -289 2092 -284
rect 1580 -328 1585 -323
rect 1595 -328 1600 -323
rect 1723 -306 1728 -301
rect 1757 -306 1762 -301
rect 2215 -311 2220 -306
rect 2230 -311 2235 -306
rect 2127 -434 2132 -429
rect 2161 -434 2166 -429
rect 1989 -452 1994 -447
rect 2004 -452 2009 -447
rect 2044 -473 2049 -468
rect 2078 -473 2083 -468
rect 2206 -495 2211 -490
rect 2221 -495 2226 -490
<< pdcontact >>
rect 929 1057 934 1062
rect 947 1057 952 1062
rect 966 1057 971 1062
rect 870 1042 875 1047
rect 885 1042 890 1047
rect 661 956 666 961
rect 725 956 730 961
rect 771 960 776 965
rect 786 960 791 965
rect 828 961 833 966
rect 843 961 848 966
rect 627 757 632 762
rect 642 757 647 762
rect 682 753 687 758
rect 698 753 703 758
rect 714 753 719 758
rect 730 753 735 758
rect 746 753 751 758
rect 762 753 767 758
rect 816 757 821 762
rect 831 757 836 762
rect 205 721 210 726
rect 220 721 225 726
rect 264 721 269 726
rect 279 721 284 726
rect 875 753 880 758
rect 891 753 896 758
rect 907 753 912 758
rect 923 753 928 758
rect 939 753 944 758
rect 974 757 979 762
rect 989 757 994 762
rect 1037 752 1042 757
rect 1053 752 1058 757
rect 1069 752 1074 757
rect 1085 752 1090 757
rect 1191 754 1196 759
rect 1209 754 1214 759
rect 1228 754 1233 759
rect 315 717 320 722
rect 349 717 354 722
rect 1132 739 1137 744
rect 1147 739 1152 744
rect 1865 728 1870 733
rect 1884 728 1889 733
rect 1902 728 1907 733
rect 2001 728 2006 733
rect 2020 728 2025 733
rect 2038 728 2043 733
rect 2147 730 2152 735
rect 2166 730 2171 735
rect 2184 730 2189 735
rect 2294 730 2299 735
rect 2313 730 2318 735
rect 2331 730 2336 735
rect 1946 713 1951 718
rect 1961 713 1966 718
rect 2082 713 2087 718
rect 2097 713 2102 718
rect 2228 715 2233 720
rect 2243 715 2248 720
rect 2506 729 2511 734
rect 2525 729 2530 734
rect 2543 729 2548 734
rect 2642 729 2647 734
rect 2661 729 2666 734
rect 2679 729 2684 734
rect 2788 731 2793 736
rect 2807 731 2812 736
rect 2825 731 2830 736
rect 2935 731 2940 736
rect 2954 731 2959 736
rect 2972 731 2977 736
rect 2375 715 2380 720
rect 2390 715 2395 720
rect 398 678 403 683
rect 432 678 437 683
rect 477 678 482 683
rect 492 678 497 683
rect 2587 714 2592 719
rect 2602 714 2607 719
rect 2723 714 2728 719
rect 2738 714 2743 719
rect 2869 716 2874 721
rect 2884 716 2889 721
rect 3016 716 3021 721
rect 3031 716 3036 721
rect 1865 620 1870 625
rect 1884 620 1889 625
rect 1902 620 1907 625
rect 2009 620 2014 625
rect 2028 620 2033 625
rect 2046 620 2051 625
rect 2158 622 2163 627
rect 2177 622 2182 627
rect 2195 622 2200 627
rect 2303 623 2308 628
rect 2322 623 2327 628
rect 2340 623 2345 628
rect 1946 605 1951 610
rect 1961 605 1966 610
rect 2090 605 2095 610
rect 2105 605 2110 610
rect 2239 607 2244 612
rect 2254 607 2259 612
rect 2384 608 2389 613
rect 2399 608 2404 613
rect 1558 550 1563 555
rect 1577 550 1582 555
rect 1595 550 1600 555
rect 202 499 207 504
rect 217 499 222 504
rect 261 499 266 504
rect 276 499 281 504
rect 1637 536 1642 541
rect 1652 536 1657 541
rect 744 508 749 513
rect 762 508 767 513
rect 781 508 786 513
rect 891 508 896 513
rect 909 508 914 513
rect 928 508 933 513
rect 312 495 317 500
rect 346 495 351 500
rect 685 493 690 498
rect 700 493 705 498
rect 832 493 837 498
rect 847 493 852 498
rect 1037 506 1042 511
rect 1055 506 1060 511
rect 1074 506 1079 511
rect 1173 506 1178 511
rect 1191 506 1196 511
rect 1210 506 1215 511
rect 978 491 983 496
rect 993 491 998 496
rect 395 456 400 461
rect 429 456 434 461
rect 474 456 479 461
rect 489 456 494 461
rect 1114 491 1119 496
rect 1129 491 1134 496
rect 2266 440 2271 445
rect 2285 440 2290 445
rect 2303 440 2308 445
rect 2402 440 2407 445
rect 2421 440 2426 445
rect 2439 440 2444 445
rect 2548 442 2553 447
rect 2567 442 2572 447
rect 2585 442 2590 447
rect 2695 442 2700 447
rect 2714 442 2719 447
rect 2732 442 2737 447
rect 1557 432 1562 437
rect 1576 432 1581 437
rect 1594 432 1599 437
rect 735 401 740 406
rect 753 401 758 406
rect 772 401 777 406
rect 676 386 681 391
rect 691 386 696 391
rect 880 400 885 405
rect 898 400 903 405
rect 917 400 922 405
rect 1636 417 1641 422
rect 1651 417 1656 422
rect 2347 425 2352 430
rect 2362 425 2367 430
rect 2483 425 2488 430
rect 2498 425 2503 430
rect 2629 427 2634 432
rect 2644 427 2649 432
rect 2776 427 2781 432
rect 2791 427 2796 432
rect 821 385 826 390
rect 836 385 841 390
rect 1029 398 1034 403
rect 1047 398 1052 403
rect 1066 398 1071 403
rect 1173 398 1178 403
rect 1191 398 1196 403
rect 1210 398 1215 403
rect 970 383 975 388
rect 985 383 990 388
rect 1114 383 1119 388
rect 1129 383 1134 388
rect 1409 397 1414 402
rect 1424 397 1429 402
rect 1447 397 1452 402
rect 1462 397 1467 402
rect 10 326 15 331
rect 25 326 30 331
rect 2005 362 2010 367
rect 2019 362 2024 367
rect 2029 362 2034 367
rect 2043 362 2048 367
rect 2074 364 2079 369
rect 2089 364 2094 369
rect 69 322 74 327
rect 85 322 90 327
rect 101 322 106 327
rect 117 322 122 327
rect 133 322 138 327
rect 205 314 210 319
rect 220 314 225 319
rect 264 314 269 319
rect 279 314 284 319
rect 1556 328 1561 333
rect 1575 328 1580 333
rect 1593 328 1598 333
rect 2266 332 2271 337
rect 2285 332 2290 337
rect 2303 332 2308 337
rect 2410 332 2415 337
rect 2429 332 2434 337
rect 2447 332 2452 337
rect 2559 334 2564 339
rect 2578 334 2583 339
rect 2596 334 2601 339
rect 2704 335 2709 340
rect 2723 335 2728 340
rect 2741 335 2746 340
rect 315 310 320 315
rect 349 310 354 315
rect 1637 313 1642 318
rect 1652 313 1657 318
rect 2347 317 2352 322
rect 2362 317 2367 322
rect 2491 317 2496 322
rect 2506 317 2511 322
rect 2640 319 2645 324
rect 2655 319 2660 324
rect 2785 320 2790 325
rect 2800 320 2805 325
rect 398 271 403 276
rect 432 271 437 276
rect 477 271 482 276
rect 492 271 497 276
rect 1556 232 1561 237
rect 1575 232 1580 237
rect 1593 232 1598 237
rect 1636 217 1641 222
rect 1651 217 1656 222
rect 205 139 210 144
rect 220 139 225 144
rect 264 139 269 144
rect 279 139 284 144
rect 315 135 320 140
rect 349 135 354 140
rect 2016 109 2021 114
rect 2031 109 2036 114
rect 398 96 403 101
rect 432 96 437 101
rect 477 96 482 101
rect 492 96 497 101
rect 2071 105 2076 110
rect 2105 105 2110 110
rect 2154 66 2159 71
rect 2188 66 2193 71
rect 2233 66 2238 71
rect 2248 66 2253 71
rect 1468 3 1473 8
rect 1483 3 1488 8
rect 1531 -1 1536 4
rect 1579 -1 1584 4
rect 2010 -74 2015 -69
rect 2025 -74 2030 -69
rect 2065 -78 2070 -73
rect 2099 -78 2104 -73
rect 1353 -115 1358 -110
rect 1371 -115 1376 -110
rect 1390 -115 1395 -110
rect 1294 -130 1299 -125
rect 1309 -130 1314 -125
rect 1499 -117 1504 -112
rect 1517 -117 1522 -112
rect 1536 -117 1541 -112
rect 1635 -117 1640 -112
rect 1653 -117 1658 -112
rect 1672 -117 1677 -112
rect 1440 -132 1445 -127
rect 1455 -132 1460 -127
rect 1576 -132 1581 -127
rect 1591 -132 1596 -127
rect 2148 -117 2153 -112
rect 2182 -117 2187 -112
rect 2227 -117 2232 -112
rect 2242 -117 2247 -112
rect 1385 -267 1390 -262
rect 1419 -267 1424 -262
rect 1467 -263 1472 -258
rect 1482 -263 1487 -258
rect 1998 -246 2003 -241
rect 2013 -246 2018 -241
rect 2053 -250 2058 -245
rect 2087 -250 2092 -245
rect 1723 -267 1728 -262
rect 1757 -267 1762 -262
rect 1799 -263 1804 -258
rect 1814 -263 1819 -258
rect 1242 -306 1247 -301
rect 1257 -306 1262 -301
rect 1302 -306 1307 -301
rect 1336 -306 1341 -301
rect 1580 -306 1585 -301
rect 1595 -306 1600 -301
rect 1640 -306 1645 -301
rect 1674 -306 1679 -301
rect 2136 -289 2141 -284
rect 2170 -289 2175 -284
rect 2215 -289 2220 -284
rect 2230 -289 2235 -284
rect 1989 -430 1994 -425
rect 2004 -430 2009 -425
rect 2044 -434 2049 -429
rect 2078 -434 2083 -429
rect 2127 -473 2132 -468
rect 2161 -473 2166 -468
rect 2206 -473 2211 -468
rect 2221 -473 2226 -468
<< nsubstratencontact >>
rect 975 1057 980 1062
rect 897 1042 902 1047
rect 737 956 742 961
rect 759 960 764 965
rect 816 961 821 966
rect 654 757 659 762
rect 843 757 848 762
rect 193 721 198 726
rect 291 721 296 726
rect 863 753 868 758
rect 1001 757 1006 762
rect 1027 752 1032 757
rect 1237 754 1242 759
rect 303 717 308 722
rect 1159 739 1164 744
rect 1856 728 1861 733
rect 1992 728 1997 733
rect 2139 730 2143 735
rect 2285 730 2290 735
rect 1934 713 1939 718
rect 2070 713 2075 718
rect 2216 715 2221 720
rect 2497 729 2502 734
rect 2633 729 2638 734
rect 2779 731 2784 736
rect 2926 731 2931 736
rect 2363 715 2368 720
rect 383 676 389 682
rect 465 678 470 683
rect 2575 714 2580 719
rect 2711 714 2716 719
rect 2857 716 2862 721
rect 3004 716 3009 721
rect 1856 620 1861 625
rect 2000 620 2005 625
rect 2149 622 2154 627
rect 2294 623 2299 628
rect 1934 605 1939 610
rect 2078 605 2083 610
rect 2227 607 2232 612
rect 2372 608 2377 613
rect 1549 550 1554 555
rect 190 499 195 504
rect 288 499 293 504
rect 1625 536 1630 541
rect 790 508 795 513
rect 937 508 942 513
rect 300 495 305 500
rect 712 493 717 498
rect 859 493 864 498
rect 1083 506 1088 511
rect 1219 506 1224 511
rect 1005 491 1010 496
rect 380 457 386 462
rect 462 456 467 461
rect 1141 491 1146 496
rect 2257 440 2262 445
rect 2393 440 2398 445
rect 2539 442 2544 447
rect 2686 442 2691 447
rect 1548 432 1553 437
rect 781 401 786 406
rect 703 386 708 391
rect 926 400 931 405
rect 1624 417 1629 422
rect 2335 425 2340 430
rect 2471 425 2476 430
rect 2617 427 2622 432
rect 2764 427 2769 432
rect 848 385 853 390
rect 1075 398 1080 403
rect 1219 398 1224 403
rect 997 383 1002 388
rect 1141 383 1146 388
rect 1397 397 1402 402
rect 37 326 42 331
rect 1995 362 2000 367
rect 2062 364 2067 369
rect 57 322 62 327
rect 168 314 173 319
rect 291 314 296 319
rect 1547 328 1552 333
rect 2257 332 2262 337
rect 2401 332 2406 337
rect 2550 334 2555 339
rect 2695 335 2700 340
rect 303 310 308 315
rect 1625 313 1630 318
rect 2335 317 2340 322
rect 2479 317 2484 322
rect 2628 319 2633 324
rect 2773 320 2778 325
rect 383 269 388 275
rect 465 271 470 276
rect 1547 232 1552 237
rect 1624 217 1629 222
rect 193 139 198 144
rect 291 139 296 144
rect 303 135 308 140
rect 2043 109 2048 114
rect 383 96 388 101
rect 465 96 470 101
rect 2059 105 2064 110
rect 2139 64 2144 69
rect 2221 66 2226 71
rect 1495 3 1500 8
rect 1522 -1 1527 4
rect 2053 -78 2058 -73
rect 1399 -115 1404 -110
rect 1321 -130 1326 -125
rect 1545 -117 1550 -112
rect 1681 -117 1686 -112
rect 1467 -132 1472 -127
rect 1603 -132 1608 -127
rect 2133 -119 2138 -114
rect 2215 -117 2220 -112
rect 1431 -267 1436 -262
rect 1455 -263 1460 -258
rect 2041 -250 2046 -245
rect 1769 -267 1774 -262
rect 1787 -263 1792 -258
rect 1269 -306 1274 -301
rect 1351 -308 1356 -303
rect 1607 -306 1612 -301
rect 1689 -308 1694 -303
rect 2121 -291 2126 -286
rect 2203 -289 2208 -284
rect 2032 -434 2037 -429
rect 2112 -475 2117 -470
rect 2194 -473 2199 -468
<< polysilicon >>
rect 936 1062 941 1076
rect 959 1062 964 1076
rect 878 1047 883 1050
rect 878 1033 883 1042
rect 936 1033 941 1057
rect 959 1033 964 1057
rect 878 1029 882 1033
rect 878 1025 883 1029
rect 878 1015 883 1020
rect 936 1009 941 1028
rect 959 1009 964 1028
rect 778 965 783 968
rect 835 966 840 969
rect 669 961 674 964
rect 685 961 690 964
rect 701 961 706 964
rect 717 961 722 964
rect 669 925 674 956
rect 685 925 690 956
rect 701 925 706 956
rect 717 925 722 956
rect 778 951 783 960
rect 835 952 840 961
rect 779 947 783 951
rect 836 948 840 952
rect 778 943 783 947
rect 835 944 840 948
rect 778 933 783 938
rect 835 934 840 939
rect 669 909 674 920
rect 685 909 690 920
rect 701 909 706 920
rect 717 910 722 920
rect 635 762 640 765
rect 690 758 695 762
rect 706 758 711 762
rect 722 758 727 777
rect 738 758 743 777
rect 824 762 829 765
rect 754 758 759 762
rect 635 748 640 757
rect 883 758 888 777
rect 899 758 904 777
rect 915 758 920 762
rect 931 758 936 777
rect 982 762 987 765
rect 341 743 379 744
rect 635 744 639 748
rect 384 743 429 744
rect 341 739 429 743
rect 635 740 640 744
rect 212 726 217 729
rect 272 726 277 729
rect 323 722 328 726
rect 341 722 346 739
rect 406 722 411 726
rect 424 722 429 739
rect 635 730 640 735
rect 690 724 695 753
rect 706 724 711 753
rect 722 724 727 753
rect 738 724 743 753
rect 754 724 759 753
rect 824 748 829 757
rect 1045 757 1050 762
rect 1061 757 1066 779
rect 1077 757 1082 777
rect 1198 759 1203 773
rect 1221 759 1226 773
rect 824 744 828 748
rect 824 740 829 744
rect 824 730 829 735
rect 883 724 888 753
rect 899 724 904 753
rect 915 724 920 753
rect 931 724 936 753
rect 982 748 987 757
rect 982 744 986 748
rect 982 740 987 744
rect 982 730 987 735
rect 212 712 217 721
rect 213 708 217 712
rect 212 704 217 708
rect 272 712 277 721
rect 1045 723 1050 752
rect 1061 723 1066 752
rect 1077 723 1082 752
rect 1140 744 1145 747
rect 1140 730 1145 739
rect 1198 730 1203 754
rect 1221 730 1226 754
rect 1872 733 1877 747
rect 1895 733 1900 747
rect 2008 733 2013 747
rect 2031 733 2036 747
rect 2154 735 2159 749
rect 2177 735 2182 749
rect 2301 735 2306 749
rect 2324 735 2329 749
rect 1140 726 1144 730
rect 272 708 276 712
rect 272 704 277 708
rect 323 705 328 717
rect 341 713 346 717
rect 406 705 411 717
rect 424 713 429 717
rect 324 700 346 705
rect 406 700 429 705
rect 690 700 695 719
rect 212 694 217 699
rect 272 694 277 699
rect 304 688 328 693
rect 304 680 309 688
rect 323 683 328 688
rect 341 683 346 700
rect 406 683 411 687
rect 424 683 429 700
rect 706 699 711 719
rect 722 702 727 719
rect 738 702 743 719
rect 754 699 759 719
rect 883 712 888 719
rect 899 712 904 719
rect 915 702 920 719
rect 931 702 936 719
rect 1140 722 1145 726
rect 2513 734 2518 748
rect 2536 734 2541 748
rect 2649 734 2654 748
rect 2672 734 2677 748
rect 2795 736 2800 750
rect 2818 736 2823 750
rect 2942 736 2947 750
rect 2965 736 2970 750
rect 1045 703 1050 718
rect 1061 704 1066 718
rect 1077 704 1082 718
rect 1140 712 1145 717
rect 1198 706 1203 725
rect 1221 706 1226 725
rect 1872 704 1877 728
rect 1895 704 1900 728
rect 1953 718 1958 721
rect 1953 704 1958 713
rect 2008 704 2013 728
rect 2031 704 2036 728
rect 2089 718 2094 721
rect 2089 704 2094 713
rect 2154 706 2159 730
rect 2177 706 2182 730
rect 2235 720 2240 723
rect 2235 706 2240 715
rect 2301 706 2306 730
rect 2324 706 2329 730
rect 2382 720 2387 723
rect 2382 706 2387 715
rect 1954 700 1958 704
rect 484 683 489 686
rect 323 660 328 678
rect 341 672 346 678
rect 1872 680 1877 699
rect 406 660 411 678
rect 323 655 411 660
rect 424 643 429 678
rect 484 669 489 678
rect 1895 680 1900 699
rect 1953 696 1958 700
rect 2090 700 2094 704
rect 2236 702 2240 706
rect 1953 686 1958 691
rect 2008 680 2013 699
rect 2031 680 2036 699
rect 2089 696 2094 700
rect 2089 686 2094 691
rect 2154 682 2159 701
rect 2177 682 2182 701
rect 2235 698 2240 702
rect 2383 702 2387 706
rect 2513 705 2518 729
rect 2536 705 2541 729
rect 2594 719 2599 722
rect 2594 705 2599 714
rect 2649 705 2654 729
rect 2672 705 2677 729
rect 2730 719 2735 722
rect 2730 705 2735 714
rect 2795 707 2800 731
rect 2818 707 2823 731
rect 2876 721 2881 724
rect 2876 707 2881 716
rect 2942 707 2947 731
rect 2965 707 2970 731
rect 3023 721 3028 724
rect 3023 707 3028 716
rect 2235 688 2240 693
rect 2301 682 2306 701
rect 2324 682 2329 701
rect 2382 698 2387 702
rect 2595 701 2599 705
rect 2382 688 2387 693
rect 2513 681 2518 700
rect 2536 681 2541 700
rect 2594 697 2599 701
rect 2731 701 2735 705
rect 2877 703 2881 707
rect 2594 687 2599 692
rect 2649 681 2654 700
rect 2672 681 2677 700
rect 2730 697 2735 701
rect 2730 687 2735 692
rect 2795 683 2800 702
rect 2818 683 2823 702
rect 2876 699 2881 703
rect 3024 703 3028 707
rect 2876 689 2881 694
rect 2942 683 2947 702
rect 2965 683 2970 702
rect 3023 699 3028 703
rect 3023 689 3028 694
rect 485 665 489 669
rect 484 661 489 665
rect 484 651 489 656
rect 1872 625 1877 639
rect 1895 625 1900 639
rect 2016 625 2021 639
rect 2039 625 2044 639
rect 2165 627 2170 641
rect 2188 627 2193 641
rect 2310 628 2315 642
rect 2333 628 2338 642
rect 1872 596 1877 620
rect 1895 596 1900 620
rect 1953 610 1958 613
rect 1953 596 1958 605
rect 2016 596 2021 620
rect 2039 596 2044 620
rect 2097 610 2102 613
rect 2097 596 2102 605
rect 2165 598 2170 622
rect 2188 598 2193 622
rect 2246 612 2251 615
rect 2246 598 2251 607
rect 2310 599 2315 623
rect 2333 599 2338 623
rect 2391 613 2396 616
rect 2391 599 2396 608
rect 1954 592 1958 596
rect 1872 572 1877 591
rect 1565 555 1570 569
rect 1588 555 1593 569
rect 1895 572 1900 591
rect 1953 588 1958 592
rect 2098 592 2102 596
rect 2247 594 2251 598
rect 2392 595 2396 599
rect 1953 578 1958 583
rect 2016 572 2021 591
rect 2039 572 2044 591
rect 2097 588 2102 592
rect 2097 578 2102 583
rect 2165 574 2170 593
rect 2188 574 2193 593
rect 2246 590 2251 594
rect 2246 580 2251 585
rect 2310 575 2315 594
rect 2333 575 2338 594
rect 2391 591 2396 595
rect 2391 581 2396 586
rect 338 521 376 522
rect 381 521 426 522
rect 338 517 426 521
rect 209 504 214 507
rect 269 504 274 507
rect 320 500 325 504
rect 338 500 343 517
rect 403 500 408 504
rect 421 500 426 517
rect 751 513 756 527
rect 774 513 779 527
rect 898 513 903 527
rect 921 513 926 527
rect 1565 526 1570 550
rect 1588 526 1593 550
rect 1644 541 1649 544
rect 1644 527 1649 536
rect 1044 511 1049 525
rect 1067 511 1072 525
rect 1180 511 1185 525
rect 1203 511 1208 525
rect 1645 523 1649 527
rect 209 490 214 499
rect 210 486 214 490
rect 209 482 214 486
rect 269 490 274 499
rect 693 498 698 501
rect 269 486 273 490
rect 269 482 274 486
rect 320 483 325 495
rect 338 491 343 495
rect 403 483 408 495
rect 421 491 426 495
rect 693 484 698 493
rect 751 484 756 508
rect 774 484 779 508
rect 840 498 845 501
rect 840 484 845 493
rect 898 484 903 508
rect 921 484 926 508
rect 986 496 991 499
rect 321 478 343 483
rect 403 478 426 483
rect 209 472 214 477
rect 269 472 274 477
rect 301 466 325 471
rect 301 458 306 466
rect 320 461 325 466
rect 338 461 343 478
rect 403 461 408 465
rect 421 461 426 478
rect 693 480 697 484
rect 693 476 698 480
rect 840 480 844 484
rect 693 466 698 471
rect 481 461 486 464
rect 751 460 756 479
rect 320 438 325 456
rect 338 450 343 456
rect 403 438 408 456
rect 320 433 408 438
rect 421 421 426 456
rect 481 447 486 456
rect 774 460 779 479
rect 840 476 845 480
rect 986 482 991 491
rect 1044 482 1049 506
rect 1067 482 1072 506
rect 1122 496 1127 499
rect 1122 482 1127 491
rect 1180 482 1185 506
rect 1203 482 1208 506
rect 1565 502 1570 521
rect 1588 502 1593 521
rect 1644 519 1649 523
rect 1644 510 1649 514
rect 840 466 845 471
rect 898 460 903 479
rect 921 460 926 479
rect 986 478 990 482
rect 986 474 991 478
rect 1122 478 1126 482
rect 986 464 991 469
rect 1044 458 1049 477
rect 1067 458 1072 477
rect 1122 474 1127 478
rect 1122 464 1127 469
rect 1180 458 1185 477
rect 1203 458 1208 477
rect 482 443 486 447
rect 481 439 486 443
rect 1564 437 1569 451
rect 1587 437 1592 451
rect 2273 445 2278 459
rect 2296 445 2301 459
rect 2409 445 2414 459
rect 2432 445 2437 459
rect 2555 447 2560 461
rect 2578 447 2583 461
rect 2702 447 2707 461
rect 2725 447 2730 461
rect 481 429 486 434
rect 742 406 747 420
rect 765 406 770 420
rect 887 405 892 419
rect 910 405 915 419
rect 684 391 689 394
rect 684 377 689 386
rect 742 377 747 401
rect 765 377 770 401
rect 1036 403 1041 417
rect 1059 403 1064 417
rect 1180 403 1185 417
rect 1203 403 1208 417
rect 1564 408 1569 432
rect 1587 408 1592 432
rect 1643 422 1648 425
rect 1643 408 1648 417
rect 2273 416 2278 440
rect 2296 416 2301 440
rect 2354 430 2359 433
rect 2354 416 2359 425
rect 2409 416 2414 440
rect 2432 416 2437 440
rect 2490 430 2495 433
rect 2490 416 2495 425
rect 2555 418 2560 442
rect 2578 418 2583 442
rect 2636 432 2641 435
rect 2636 418 2641 427
rect 2702 418 2707 442
rect 2725 418 2730 442
rect 2783 432 2788 435
rect 2783 418 2788 427
rect 2355 412 2359 416
rect 829 390 834 393
rect 684 373 688 377
rect 684 369 689 373
rect 829 376 834 385
rect 887 376 892 400
rect 910 376 915 400
rect 1416 402 1421 405
rect 1454 402 1459 405
rect 1644 404 1648 408
rect 978 388 983 391
rect 829 372 833 376
rect 684 359 689 364
rect 742 353 747 372
rect 765 353 770 372
rect 829 368 834 372
rect 978 374 983 383
rect 1036 374 1041 398
rect 1059 374 1064 398
rect 1122 388 1127 391
rect 1122 374 1127 383
rect 1180 374 1185 398
rect 1203 374 1208 398
rect 1416 388 1421 397
rect 1454 388 1459 397
rect 1417 384 1421 388
rect 1455 384 1459 388
rect 1416 380 1421 384
rect 1454 380 1459 384
rect 1564 384 1569 403
rect 1587 384 1592 403
rect 1643 400 1648 404
rect 1643 390 1648 395
rect 829 358 834 363
rect 887 352 892 371
rect 910 352 915 371
rect 978 370 982 374
rect 978 366 983 370
rect 1122 370 1126 374
rect 978 356 983 361
rect 1036 350 1041 369
rect 18 331 23 334
rect 77 327 82 346
rect 93 327 98 346
rect 1059 350 1064 369
rect 1122 366 1127 370
rect 1416 370 1421 375
rect 1454 370 1459 375
rect 1122 356 1127 361
rect 1180 350 1185 369
rect 1203 350 1208 369
rect 2012 367 2017 375
rect 2036 367 2041 401
rect 2273 392 2278 411
rect 2296 392 2301 411
rect 2354 408 2359 412
rect 2491 412 2495 416
rect 2637 414 2641 418
rect 2354 398 2359 403
rect 2409 392 2414 411
rect 2432 392 2437 411
rect 2490 408 2495 412
rect 2490 398 2495 403
rect 2555 394 2560 413
rect 2578 394 2583 413
rect 2636 410 2641 414
rect 2784 414 2788 418
rect 2636 400 2641 405
rect 2702 394 2707 413
rect 2725 394 2730 413
rect 2783 410 2788 414
rect 2783 400 2788 405
rect 2081 369 2086 372
rect 2012 352 2017 362
rect 2013 347 2017 352
rect 341 336 379 337
rect 384 336 429 337
rect 341 332 429 336
rect 1563 333 1568 347
rect 1586 333 1591 347
rect 109 327 114 331
rect 125 327 130 331
rect 18 317 23 326
rect 18 313 22 317
rect 18 309 23 313
rect 18 299 23 304
rect 77 293 82 322
rect 93 293 98 322
rect 109 293 114 322
rect 125 293 130 322
rect 212 319 217 322
rect 272 319 277 322
rect 323 315 328 319
rect 341 315 346 332
rect 406 315 411 319
rect 424 315 429 332
rect 2012 330 2017 347
rect 2036 330 2041 362
rect 2081 355 2086 364
rect 2082 351 2086 355
rect 2081 347 2086 351
rect 2081 337 2086 342
rect 2273 337 2278 351
rect 2296 337 2301 351
rect 2417 337 2422 351
rect 2440 337 2445 351
rect 2566 339 2571 353
rect 2589 339 2594 353
rect 2711 340 2716 354
rect 2734 340 2739 354
rect 212 305 217 314
rect 213 301 217 305
rect 212 297 217 301
rect 272 305 277 314
rect 272 301 276 305
rect 272 297 277 301
rect 323 298 328 310
rect 341 306 346 310
rect 406 298 411 310
rect 424 306 429 310
rect 1563 304 1568 328
rect 1586 304 1591 328
rect 2012 321 2017 325
rect 2036 321 2041 325
rect 1644 318 1649 321
rect 1644 304 1649 313
rect 2273 308 2278 332
rect 2296 308 2301 332
rect 2354 322 2359 325
rect 2354 308 2359 317
rect 2417 308 2422 332
rect 2440 308 2445 332
rect 2498 322 2503 325
rect 2498 308 2503 317
rect 2566 310 2571 334
rect 2589 310 2594 334
rect 2647 324 2652 327
rect 2647 310 2652 319
rect 2711 311 2716 335
rect 2734 311 2739 335
rect 2792 325 2797 328
rect 2792 311 2797 320
rect 1645 300 1649 304
rect 2355 304 2359 308
rect 324 293 346 298
rect 406 293 429 298
rect 77 281 82 288
rect 93 281 98 288
rect 109 271 114 288
rect 125 271 130 288
rect 212 287 217 292
rect 272 287 277 292
rect 304 281 328 286
rect 304 273 309 281
rect 323 276 328 281
rect 341 276 346 293
rect 406 276 411 280
rect 424 276 429 293
rect 1563 280 1568 299
rect 484 276 489 279
rect 323 253 328 271
rect 341 265 346 271
rect 1586 280 1591 299
rect 1644 296 1649 300
rect 1644 286 1649 291
rect 2273 284 2278 303
rect 2296 284 2301 303
rect 2354 300 2359 304
rect 2499 304 2503 308
rect 2648 306 2652 310
rect 2793 307 2797 311
rect 2354 290 2359 295
rect 2417 284 2422 303
rect 2440 284 2445 303
rect 2498 300 2503 304
rect 2498 290 2503 295
rect 2566 286 2571 305
rect 2589 286 2594 305
rect 2647 302 2652 306
rect 2647 292 2652 297
rect 2711 287 2716 306
rect 2734 287 2739 306
rect 2792 303 2797 307
rect 2792 293 2797 298
rect 406 253 411 271
rect 323 248 411 253
rect 424 236 429 271
rect 484 262 489 271
rect 485 258 489 262
rect 484 254 489 258
rect 484 244 489 249
rect 1563 237 1568 251
rect 1586 237 1591 251
rect 1563 208 1568 232
rect 1586 208 1591 232
rect 1643 222 1648 225
rect 1643 208 1648 217
rect 1644 204 1648 208
rect 1563 184 1568 203
rect 1586 184 1591 203
rect 1643 200 1648 204
rect 1643 190 1648 195
rect 341 161 379 162
rect 384 161 429 162
rect 341 157 429 161
rect 212 144 217 147
rect 272 144 277 147
rect 323 140 328 144
rect 341 140 346 157
rect 406 140 411 144
rect 424 140 429 157
rect 212 130 217 139
rect 213 126 217 130
rect 212 122 217 126
rect 272 130 277 139
rect 272 126 276 130
rect 272 122 277 126
rect 323 123 328 135
rect 341 131 346 135
rect 406 123 411 135
rect 424 131 429 135
rect 2097 131 2135 132
rect 2140 131 2185 132
rect 2097 127 2185 131
rect 324 118 346 123
rect 406 118 429 123
rect 212 112 217 117
rect 272 112 277 117
rect 304 106 328 111
rect 304 98 309 106
rect 323 101 328 106
rect 341 101 346 118
rect 406 101 411 105
rect 424 101 429 118
rect 2024 114 2029 117
rect 2079 110 2084 114
rect 2097 110 2102 127
rect 2162 110 2167 114
rect 2180 110 2185 127
rect 484 101 489 104
rect 2024 100 2029 109
rect 2024 96 2028 100
rect 323 78 328 96
rect 341 90 346 96
rect 406 78 411 96
rect 323 73 411 78
rect 424 61 429 96
rect 484 87 489 96
rect 2024 92 2029 96
rect 2079 93 2084 105
rect 2097 101 2102 105
rect 2162 93 2167 105
rect 2180 101 2185 105
rect 2080 88 2102 93
rect 2162 88 2185 93
rect 485 83 489 87
rect 484 79 489 83
rect 2024 82 2029 87
rect 2060 76 2084 81
rect 484 69 489 74
rect 2060 68 2065 76
rect 2079 71 2084 76
rect 2097 71 2102 88
rect 2162 71 2167 75
rect 2180 71 2185 88
rect 2240 71 2245 74
rect 2079 48 2084 66
rect 2097 60 2102 66
rect 2162 48 2167 66
rect 2079 43 2167 48
rect 2180 31 2185 66
rect 2240 57 2245 66
rect 2241 53 2245 57
rect 2240 49 2245 53
rect 2240 39 2245 44
rect 1476 8 1481 11
rect 1539 4 1544 7
rect 1555 4 1560 7
rect 1571 4 1576 7
rect 1476 -6 1481 3
rect 1476 -10 1480 -6
rect 1476 -14 1481 -10
rect 1476 -24 1481 -19
rect 1539 -32 1544 -1
rect 1555 -32 1560 -1
rect 1571 -32 1576 -1
rect 1539 -48 1544 -37
rect 1555 -48 1560 -37
rect 1571 -48 1576 -37
rect 2091 -52 2129 -51
rect 2134 -52 2179 -51
rect 2091 -56 2179 -52
rect 2018 -69 2023 -66
rect 2073 -73 2078 -69
rect 2091 -73 2096 -56
rect 2156 -73 2161 -69
rect 2174 -73 2179 -56
rect 2018 -83 2023 -74
rect 2018 -87 2022 -83
rect 2018 -91 2023 -87
rect 2073 -90 2078 -78
rect 2091 -82 2096 -78
rect 2156 -90 2161 -78
rect 2174 -82 2179 -78
rect 2074 -95 2096 -90
rect 2156 -95 2179 -90
rect 1360 -110 1365 -96
rect 1383 -110 1388 -96
rect 1506 -112 1511 -98
rect 1529 -112 1534 -98
rect 1642 -112 1647 -98
rect 1665 -112 1670 -98
rect 2018 -101 2023 -96
rect 2054 -107 2078 -102
rect 1302 -125 1307 -122
rect 1302 -139 1307 -130
rect 1360 -139 1365 -115
rect 1383 -139 1388 -115
rect 2054 -115 2059 -107
rect 2073 -112 2078 -107
rect 2091 -112 2096 -95
rect 2156 -112 2161 -108
rect 2174 -112 2179 -95
rect 2234 -112 2239 -109
rect 1448 -127 1453 -124
rect 1302 -143 1306 -139
rect 1302 -147 1307 -143
rect 1448 -141 1453 -132
rect 1506 -141 1511 -117
rect 1529 -141 1534 -117
rect 1584 -127 1589 -124
rect 1584 -141 1589 -132
rect 1642 -141 1647 -117
rect 1665 -141 1670 -117
rect 2073 -135 2078 -117
rect 2091 -123 2096 -117
rect 2156 -135 2161 -117
rect 2073 -140 2161 -135
rect 1302 -157 1307 -152
rect 1360 -163 1365 -144
rect 1383 -163 1388 -144
rect 1448 -145 1452 -141
rect 1448 -149 1453 -145
rect 1584 -145 1588 -141
rect 1448 -159 1453 -154
rect 1506 -165 1511 -146
rect 1529 -165 1534 -146
rect 1584 -149 1589 -145
rect 1584 -159 1589 -154
rect 1642 -165 1647 -146
rect 1665 -165 1670 -146
rect 2174 -152 2179 -117
rect 2234 -126 2239 -117
rect 2235 -130 2239 -126
rect 2234 -134 2239 -130
rect 2234 -144 2239 -139
rect 2079 -224 2117 -223
rect 2122 -224 2167 -223
rect 2079 -228 2167 -224
rect 1310 -241 1355 -240
rect 1360 -241 1398 -240
rect 1310 -245 1398 -241
rect 1310 -262 1315 -245
rect 1328 -262 1333 -258
rect 1393 -262 1398 -245
rect 1648 -241 1693 -240
rect 1698 -241 1736 -240
rect 2006 -241 2011 -238
rect 1648 -245 1736 -241
rect 1474 -258 1479 -255
rect 1411 -262 1416 -258
rect 1648 -262 1653 -245
rect 1666 -262 1671 -258
rect 1731 -262 1736 -245
rect 2061 -245 2066 -241
rect 2079 -245 2084 -228
rect 2144 -245 2149 -241
rect 2162 -245 2167 -228
rect 2006 -255 2011 -246
rect 1806 -258 1811 -255
rect 1749 -262 1754 -258
rect 1310 -271 1315 -267
rect 1328 -279 1333 -267
rect 1393 -271 1398 -267
rect 1411 -279 1416 -267
rect 1474 -272 1479 -263
rect 2006 -259 2010 -255
rect 2006 -263 2011 -259
rect 2061 -262 2066 -250
rect 2079 -254 2084 -250
rect 2144 -262 2149 -250
rect 2162 -254 2167 -250
rect 1648 -271 1653 -267
rect 1475 -276 1479 -272
rect 1310 -284 1333 -279
rect 1393 -284 1415 -279
rect 1474 -280 1479 -276
rect 1666 -279 1671 -267
rect 1731 -271 1736 -267
rect 1749 -279 1754 -267
rect 1806 -272 1811 -263
rect 2062 -267 2084 -262
rect 2144 -267 2167 -262
rect 1807 -276 1811 -272
rect 2006 -273 2011 -268
rect 1250 -301 1255 -298
rect 1310 -301 1315 -284
rect 1328 -301 1333 -297
rect 1393 -301 1398 -284
rect 1648 -284 1671 -279
rect 1731 -284 1753 -279
rect 1806 -280 1811 -276
rect 2042 -279 2066 -274
rect 1474 -290 1479 -285
rect 1411 -296 1435 -291
rect 1411 -301 1416 -296
rect 1250 -315 1255 -306
rect 1250 -319 1254 -315
rect 1250 -323 1255 -319
rect 1250 -333 1255 -328
rect 1310 -341 1315 -306
rect 1328 -324 1333 -306
rect 1430 -304 1435 -296
rect 1588 -301 1593 -298
rect 1648 -301 1653 -284
rect 1666 -301 1671 -297
rect 1731 -301 1736 -284
rect 1806 -290 1811 -285
rect 2042 -287 2047 -279
rect 2061 -284 2066 -279
rect 2079 -284 2084 -267
rect 2144 -284 2149 -280
rect 2162 -284 2167 -267
rect 2222 -284 2227 -281
rect 1749 -296 1773 -291
rect 1749 -301 1754 -296
rect 1393 -312 1398 -306
rect 1411 -324 1416 -306
rect 1588 -315 1593 -306
rect 1588 -319 1592 -315
rect 1588 -323 1593 -319
rect 1328 -329 1416 -324
rect 1588 -333 1593 -328
rect 1648 -341 1653 -306
rect 1666 -324 1671 -306
rect 1768 -304 1773 -296
rect 1731 -312 1736 -306
rect 1749 -324 1754 -306
rect 2061 -307 2066 -289
rect 2079 -295 2084 -289
rect 2144 -307 2149 -289
rect 2061 -312 2149 -307
rect 1666 -329 1754 -324
rect 2162 -324 2167 -289
rect 2222 -298 2227 -289
rect 2223 -302 2227 -298
rect 2222 -306 2227 -302
rect 2222 -316 2227 -311
rect 2070 -408 2108 -407
rect 2113 -408 2158 -407
rect 2070 -412 2158 -408
rect 1997 -425 2002 -422
rect 2052 -429 2057 -425
rect 2070 -429 2075 -412
rect 2135 -429 2140 -425
rect 2153 -429 2158 -412
rect 1997 -439 2002 -430
rect 1997 -443 2001 -439
rect 1997 -447 2002 -443
rect 2052 -446 2057 -434
rect 2070 -438 2075 -434
rect 2135 -446 2140 -434
rect 2153 -438 2158 -434
rect 2053 -451 2075 -446
rect 2135 -451 2158 -446
rect 1997 -457 2002 -452
rect 2033 -463 2057 -458
rect 2033 -471 2038 -463
rect 2052 -468 2057 -463
rect 2070 -468 2075 -451
rect 2135 -468 2140 -464
rect 2153 -468 2158 -451
rect 2213 -468 2218 -465
rect 2052 -491 2057 -473
rect 2070 -479 2075 -473
rect 2135 -491 2140 -473
rect 2052 -496 2140 -491
rect 2153 -508 2158 -473
rect 2213 -482 2218 -473
rect 2214 -486 2218 -482
rect 2213 -490 2218 -486
rect 2213 -500 2218 -495
<< polycontact >>
rect 882 1029 887 1033
rect 936 1003 941 1009
rect 959 1003 964 1009
rect 774 947 779 951
rect 831 948 836 952
rect 669 902 674 909
rect 685 902 690 909
rect 701 902 706 909
rect 717 903 722 910
rect 722 777 727 782
rect 738 777 744 783
rect 883 777 889 784
rect 899 777 905 784
rect 931 777 937 783
rect 1060 779 1067 785
rect 379 743 384 748
rect 639 744 644 748
rect 1075 777 1085 785
rect 828 744 833 748
rect 986 744 991 748
rect 208 708 213 712
rect 1144 726 1149 730
rect 276 708 281 712
rect 319 700 324 705
rect 915 696 922 702
rect 1043 696 1051 703
rect 1198 700 1203 706
rect 1221 700 1226 706
rect 1949 700 1954 704
rect 304 675 309 680
rect 1872 674 1877 680
rect 2085 700 2090 704
rect 2231 702 2236 706
rect 1895 674 1900 680
rect 2008 674 2013 680
rect 2031 674 2036 680
rect 2154 676 2159 682
rect 2378 702 2383 706
rect 2177 676 2182 682
rect 2301 676 2306 682
rect 2590 701 2595 705
rect 2324 676 2329 682
rect 2513 675 2518 681
rect 2726 701 2731 705
rect 2872 703 2877 707
rect 2536 675 2541 681
rect 2649 675 2654 681
rect 2672 675 2677 681
rect 2795 677 2800 683
rect 3019 703 3024 707
rect 2818 677 2823 683
rect 2942 677 2947 683
rect 2965 677 2970 683
rect 480 665 485 669
rect 424 638 429 643
rect 1949 592 1954 596
rect 1872 566 1877 572
rect 2093 592 2098 596
rect 2242 594 2247 598
rect 2387 595 2392 599
rect 1895 566 1900 572
rect 2016 566 2021 572
rect 2039 566 2044 572
rect 2165 568 2170 574
rect 2188 568 2193 574
rect 2310 569 2315 575
rect 2333 569 2338 575
rect 376 521 381 526
rect 1640 523 1645 527
rect 205 486 210 490
rect 273 486 278 490
rect 316 478 321 483
rect 301 453 306 458
rect 697 480 702 484
rect 844 480 849 484
rect 751 454 756 460
rect 1565 496 1570 502
rect 1588 496 1593 502
rect 774 454 779 460
rect 898 454 903 460
rect 990 478 995 482
rect 1126 478 1131 482
rect 921 454 926 460
rect 1044 452 1049 458
rect 1067 452 1072 458
rect 1180 452 1185 458
rect 1203 452 1208 458
rect 477 443 482 447
rect 421 416 426 421
rect 2350 412 2355 416
rect 688 373 693 377
rect 1639 404 1644 408
rect 833 372 838 376
rect 77 346 83 353
rect 93 346 99 353
rect 742 347 747 353
rect 1412 384 1417 388
rect 1450 384 1455 388
rect 1564 378 1569 384
rect 2036 401 2042 407
rect 1587 378 1592 384
rect 765 347 770 353
rect 887 346 892 352
rect 982 370 987 374
rect 1126 370 1131 374
rect 910 346 915 352
rect 1036 344 1041 350
rect 1059 344 1064 350
rect 1180 344 1185 350
rect 2273 386 2278 392
rect 2486 412 2491 416
rect 2632 414 2637 418
rect 2296 386 2301 392
rect 2409 386 2414 392
rect 2432 386 2437 392
rect 2555 388 2560 394
rect 2779 414 2784 418
rect 2578 388 2583 394
rect 2702 388 2707 394
rect 2725 388 2730 394
rect 1203 344 1208 350
rect 2008 347 2013 352
rect 379 336 384 341
rect 22 313 27 317
rect 2077 351 2082 355
rect 208 301 213 305
rect 276 301 281 305
rect 1640 300 1645 304
rect 2350 304 2355 308
rect 319 293 324 298
rect 109 265 116 271
rect 125 265 132 271
rect 304 268 309 273
rect 1563 274 1568 280
rect 1586 274 1591 280
rect 2273 278 2278 284
rect 2494 304 2499 308
rect 2643 306 2648 310
rect 2788 307 2793 311
rect 2296 278 2301 284
rect 2417 278 2422 284
rect 2440 278 2445 284
rect 2566 280 2571 286
rect 2589 280 2594 286
rect 2711 281 2716 287
rect 2734 281 2739 287
rect 480 258 485 262
rect 424 231 429 236
rect 1639 204 1644 208
rect 1563 178 1568 184
rect 1586 178 1591 184
rect 379 161 384 166
rect 208 126 213 130
rect 276 126 281 130
rect 2135 131 2140 136
rect 319 118 324 123
rect 304 93 309 98
rect 2028 96 2033 100
rect 2075 88 2080 93
rect 480 83 485 87
rect 2060 63 2065 68
rect 424 56 429 61
rect 2236 53 2241 57
rect 2180 26 2185 31
rect 1480 -10 1485 -6
rect 1539 -55 1544 -48
rect 1555 -55 1560 -48
rect 1571 -55 1576 -48
rect 2129 -52 2134 -47
rect 2022 -87 2027 -83
rect 2069 -95 2074 -90
rect 1306 -143 1311 -139
rect 2054 -120 2059 -115
rect 1360 -169 1365 -163
rect 1452 -145 1457 -141
rect 1588 -145 1593 -141
rect 1383 -169 1388 -163
rect 1506 -171 1511 -165
rect 1529 -171 1534 -165
rect 1642 -171 1647 -165
rect 2230 -130 2235 -126
rect 2174 -157 2179 -152
rect 1665 -171 1670 -165
rect 2117 -224 2122 -219
rect 1355 -241 1360 -236
rect 1693 -241 1698 -236
rect 2010 -259 2015 -255
rect 1470 -276 1475 -272
rect 1415 -284 1420 -279
rect 2057 -267 2062 -262
rect 1802 -276 1807 -272
rect 1753 -284 1758 -279
rect 1254 -319 1259 -315
rect 2042 -292 2047 -287
rect 1430 -309 1435 -304
rect 1592 -319 1597 -315
rect 1310 -346 1315 -341
rect 1768 -309 1773 -304
rect 2218 -302 2223 -298
rect 2162 -329 2167 -324
rect 1648 -346 1653 -341
rect 2108 -408 2113 -403
rect 2001 -443 2006 -439
rect 2048 -451 2053 -446
rect 2033 -476 2038 -471
rect 2209 -486 2214 -482
rect 2153 -513 2158 -508
<< metal1 >>
rect 904 1073 932 1074
rect 904 1070 990 1073
rect 904 1060 908 1070
rect 929 1069 990 1070
rect 929 1068 980 1069
rect 929 1062 934 1068
rect 966 1062 971 1068
rect 904 1059 909 1060
rect 861 1054 909 1059
rect 975 1062 980 1068
rect 885 1047 890 1054
rect 897 1047 902 1054
rect 947 1047 952 1057
rect 947 1043 957 1047
rect 870 1033 875 1042
rect 953 1039 957 1043
rect 916 1036 957 1039
rect 916 1033 919 1036
rect 953 1033 957 1036
rect 859 1029 875 1033
rect 887 1029 919 1033
rect 870 1025 875 1029
rect 927 1028 929 1031
rect 885 1016 890 1020
rect 927 1017 930 1028
rect 944 1025 947 1028
rect 971 1017 974 1031
rect 859 1011 895 1016
rect 859 1010 866 1011
rect 927 1012 974 1017
rect 859 989 864 1010
rect 936 1002 941 1003
rect 959 987 964 1003
rect 950 984 964 987
rect 809 977 857 978
rect 985 977 990 1069
rect 1247 977 1270 978
rect 647 974 1271 977
rect 647 973 1262 974
rect 647 972 800 973
rect 661 961 666 972
rect 737 961 742 972
rect 759 965 764 972
rect 771 965 776 972
rect 816 966 821 973
rect 828 966 833 973
rect 725 934 730 956
rect 786 951 791 960
rect 843 952 848 961
rect 944 952 948 960
rect 795 951 831 952
rect 756 947 774 951
rect 786 948 831 951
rect 843 948 948 952
rect 786 947 829 948
rect 756 934 759 947
rect 786 943 791 947
rect 843 944 848 948
rect 771 934 776 938
rect 828 935 833 939
rect 819 934 858 935
rect 677 930 759 934
rect 762 930 882 934
rect 677 925 682 930
rect 709 925 714 930
rect 762 929 801 930
rect 889 930 1181 934
rect 661 916 666 920
rect 693 917 698 920
rect 725 917 730 920
rect 762 917 767 929
rect 693 916 767 917
rect 661 913 767 916
rect 669 900 674 902
rect 685 898 690 902
rect 685 885 689 898
rect 701 897 706 902
rect 722 903 866 904
rect 717 899 866 903
rect 1178 903 1181 930
rect 1266 921 1271 974
rect 685 882 795 885
rect 292 873 934 875
rect 292 872 935 873
rect 292 808 295 872
rect 655 849 660 864
rect 796 849 800 864
rect 931 851 935 872
rect 141 805 295 808
rect 178 804 295 805
rect 578 837 585 840
rect 928 837 952 838
rect 578 834 1066 837
rect 94 782 186 784
rect 93 777 186 782
rect 76 354 82 763
rect 77 353 82 354
rect 93 544 99 777
rect 460 763 461 769
rect 475 763 554 769
rect 379 750 530 755
rect 178 746 372 750
rect 178 712 183 746
rect 193 734 356 738
rect 193 733 308 734
rect 193 726 198 733
rect 205 726 210 733
rect 279 726 284 733
rect 220 712 225 721
rect 291 726 296 733
rect 303 722 308 733
rect 178 709 208 712
rect 204 708 208 709
rect 220 708 229 712
rect 264 712 269 721
rect 315 722 320 734
rect 238 708 269 712
rect 281 708 287 712
rect 220 704 225 708
rect 205 695 210 699
rect 196 690 227 695
rect 238 644 242 708
rect 264 704 269 708
rect 294 708 302 712
rect 298 705 302 708
rect 349 711 354 717
rect 367 711 372 746
rect 379 748 384 750
rect 398 728 451 734
rect 398 722 403 728
rect 432 711 437 717
rect 349 706 437 711
rect 298 700 319 705
rect 279 695 284 699
rect 255 690 293 695
rect 283 653 288 690
rect 349 683 354 706
rect 304 672 309 675
rect 383 682 389 695
rect 315 653 320 678
rect 398 683 403 693
rect 432 683 437 706
rect 446 653 451 728
rect 463 690 506 695
rect 465 683 470 690
rect 477 683 482 690
rect 492 670 497 678
rect 511 670 516 750
rect 548 680 554 763
rect 578 715 585 834
rect 717 824 736 829
rect 607 698 611 823
rect 655 786 660 823
rect 717 788 725 824
rect 796 788 800 826
rect 853 794 889 801
rect 717 787 743 788
rect 717 785 744 787
rect 736 783 744 785
rect 690 777 722 782
rect 736 781 738 783
rect 882 785 888 794
rect 883 784 888 785
rect 899 784 904 789
rect 931 783 935 825
rect 1061 785 1066 834
rect 1077 803 1081 853
rect 1178 795 1182 903
rect 1265 901 1271 921
rect 1077 785 1081 792
rect 617 770 1130 774
rect 1265 772 1270 901
rect 2097 826 2104 827
rect 2097 822 2362 826
rect 2097 821 2370 822
rect 2071 802 2076 807
rect 2097 802 2104 821
rect 2071 796 2104 802
rect 1248 771 1349 772
rect 618 769 666 770
rect 642 762 647 769
rect 654 762 659 769
rect 698 758 703 770
rect 730 758 735 770
rect 762 758 767 770
rect 807 769 855 770
rect 627 748 632 757
rect 831 762 836 769
rect 682 750 687 753
rect 714 750 719 753
rect 682 749 719 750
rect 746 749 751 753
rect 622 744 632 748
rect 644 745 668 748
rect 644 744 659 745
rect 627 740 632 744
rect 642 731 647 735
rect 664 736 668 745
rect 682 745 751 749
rect 796 748 800 758
rect 843 762 848 769
rect 863 758 868 770
rect 816 748 821 757
rect 875 758 880 770
rect 907 758 912 770
rect 939 758 944 770
rect 965 769 1130 770
rect 989 762 994 769
rect 1001 762 1006 769
rect 1027 757 1032 769
rect 1053 757 1058 769
rect 1085 757 1090 769
rect 891 750 896 753
rect 876 749 896 750
rect 923 749 928 753
rect 682 736 687 745
rect 796 744 821 748
rect 833 744 852 748
rect 664 731 687 736
rect 816 740 821 744
rect 831 731 836 735
rect 848 736 852 744
rect 876 745 928 749
rect 876 736 881 745
rect 974 748 979 757
rect 1036 752 1037 757
rect 1124 756 1130 769
rect 1163 770 1194 771
rect 1241 770 1349 771
rect 1163 767 1349 770
rect 1167 756 1171 767
rect 1036 749 1042 752
rect 1069 749 1074 752
rect 1123 751 1171 756
rect 1191 765 1242 767
rect 1248 766 1349 767
rect 1191 759 1196 765
rect 1228 759 1233 765
rect 1237 759 1242 765
rect 967 744 979 748
rect 991 744 1017 748
rect 1036 744 1074 749
rect 1147 744 1152 751
rect 848 731 881 736
rect 974 740 979 744
rect 989 731 994 735
rect 1013 731 1017 744
rect 1034 731 1039 744
rect 1159 744 1164 751
rect 1209 744 1214 754
rect 1209 740 1219 744
rect 617 726 656 731
rect 651 710 656 726
rect 682 724 687 731
rect 806 726 845 731
rect 762 712 767 719
rect 840 712 845 726
rect 876 724 881 731
rect 963 726 1009 731
rect 1013 726 1039 731
rect 762 710 845 712
rect 939 717 944 719
rect 964 717 970 726
rect 939 714 970 717
rect 1005 725 1009 726
rect 939 713 949 714
rect 939 710 944 713
rect 651 707 944 710
rect 1005 711 1010 725
rect 1034 723 1039 726
rect 1132 730 1137 739
rect 1215 736 1219 740
rect 1178 733 1219 736
rect 1178 730 1181 733
rect 1215 730 1219 733
rect 1126 726 1137 730
rect 1149 726 1181 730
rect 1085 711 1090 718
rect 1132 722 1137 726
rect 1189 725 1191 728
rect 1147 713 1152 717
rect 1189 714 1192 725
rect 1206 722 1209 725
rect 1233 714 1236 728
rect 1121 711 1157 713
rect 1005 708 1157 711
rect 1005 707 1130 708
rect 1189 709 1236 714
rect 651 706 767 707
rect 840 706 944 707
rect 607 696 690 698
rect 607 694 695 696
rect 706 689 711 696
rect 754 693 759 696
rect 706 685 737 689
rect 548 678 683 680
rect 548 675 684 678
rect 477 665 480 669
rect 492 665 516 670
rect 492 661 497 665
rect 678 661 684 675
rect 728 674 736 685
rect 730 666 736 674
rect 753 680 762 693
rect 915 692 920 696
rect 1045 693 1049 696
rect 753 673 755 680
rect 728 665 736 666
rect 283 652 451 653
rect 477 652 482 656
rect 283 648 530 652
rect 446 647 530 648
rect 238 639 407 644
rect 402 634 407 639
rect 424 634 429 638
rect 402 629 429 634
rect 93 541 224 544
rect 93 540 99 541
rect 93 353 98 540
rect 507 533 514 599
rect 376 528 514 533
rect 175 524 369 528
rect 175 490 180 524
rect 190 512 353 516
rect 190 511 305 512
rect 190 504 195 511
rect 202 504 207 511
rect 276 504 281 511
rect 217 490 222 499
rect 288 504 293 511
rect 300 500 305 511
rect 175 487 205 490
rect 201 486 205 487
rect 217 486 226 490
rect 261 490 266 499
rect 312 500 317 512
rect 235 486 266 490
rect 278 488 299 490
rect 278 486 286 488
rect 217 482 222 486
rect 202 473 207 477
rect 193 468 224 473
rect 235 422 239 486
rect 261 482 266 486
rect 292 486 299 488
rect 295 483 299 486
rect 346 489 351 495
rect 364 489 369 524
rect 376 526 381 528
rect 395 506 448 512
rect 395 500 400 506
rect 429 489 434 495
rect 346 484 434 489
rect 295 478 316 483
rect 276 473 281 477
rect 252 468 290 473
rect 280 431 285 468
rect 346 461 351 484
rect 395 478 398 481
rect 388 473 403 478
rect 301 450 306 453
rect 380 462 385 473
rect 395 461 400 473
rect 429 461 434 484
rect 312 431 317 456
rect 443 431 448 506
rect 460 468 503 473
rect 462 461 467 468
rect 474 461 479 468
rect 489 448 494 456
rect 508 448 513 528
rect 474 443 477 447
rect 489 443 513 448
rect 523 465 529 647
rect 548 610 557 648
rect 677 655 684 661
rect 570 596 577 647
rect 620 623 621 630
rect 620 566 627 623
rect 552 558 628 566
rect 677 558 683 655
rect 739 617 748 642
rect 914 638 920 692
rect 1044 630 1049 693
rect 1121 685 1130 707
rect 1198 699 1203 700
rect 1221 699 1226 700
rect 1122 676 1130 685
rect 1122 675 1322 676
rect 1122 673 1325 675
rect 1318 665 1325 673
rect 739 611 1109 617
rect 789 579 815 585
rect 1102 577 1109 611
rect 727 562 958 566
rect 1319 561 1323 665
rect 676 553 683 558
rect 585 532 651 539
rect 677 510 683 553
rect 716 524 747 525
rect 794 524 894 525
rect 716 523 942 524
rect 716 522 1040 523
rect 1145 522 1176 523
rect 1343 522 1347 766
rect 1676 767 1991 771
rect 1855 766 1991 767
rect 2071 764 2076 796
rect 2097 795 2104 796
rect 2118 797 2618 802
rect 2118 777 2124 797
rect 2071 760 2132 764
rect 2188 763 2193 778
rect 2271 774 2766 780
rect 2188 760 2281 763
rect 1693 744 1700 749
rect 2827 747 2927 748
rect 2974 747 3005 748
rect 2186 746 2286 747
rect 2333 746 2364 747
rect 2779 746 3005 747
rect 2132 745 2364 746
rect 2545 745 2576 746
rect 2681 745 3005 746
rect 1904 744 1935 745
rect 2040 744 2364 745
rect 2490 744 3005 745
rect 1693 743 2830 744
rect 1693 741 2189 743
rect 1693 739 1907 741
rect 1471 566 1476 568
rect 1693 567 1700 739
rect 1835 738 1862 739
rect 1835 638 1843 738
rect 1856 733 1861 738
rect 1865 733 1870 739
rect 1902 733 1907 739
rect 1927 740 2043 741
rect 1927 730 1931 740
rect 1992 739 2043 740
rect 1992 733 1997 739
rect 1884 718 1889 728
rect 1927 725 1975 730
rect 2001 733 2006 739
rect 2038 733 2043 739
rect 2063 730 2067 741
rect 2139 735 2143 741
rect 2147 735 2152 741
rect 2184 735 2189 741
rect 2209 732 2213 743
rect 2285 741 2336 743
rect 2285 735 2290 741
rect 1879 714 1889 718
rect 1934 718 1939 725
rect 1879 710 1883 714
rect 1946 718 1951 725
rect 2020 718 2025 728
rect 2063 725 2111 730
rect 1879 707 1920 710
rect 1879 704 1883 707
rect 1917 704 1920 707
rect 1961 704 1966 713
rect 2015 714 2025 718
rect 2070 718 2075 725
rect 2015 710 2019 714
rect 2082 718 2087 725
rect 2166 720 2171 730
rect 2209 727 2257 732
rect 2294 735 2299 741
rect 2331 735 2336 741
rect 2356 742 2830 743
rect 2356 740 2548 742
rect 2356 732 2360 740
rect 2490 739 2503 740
rect 2497 734 2502 739
rect 2015 707 2056 710
rect 1862 688 1865 702
rect 1907 699 1909 702
rect 1917 700 1949 704
rect 1961 700 1980 704
rect 1889 696 1892 699
rect 1906 688 1909 699
rect 1961 696 1966 700
rect 2015 704 2019 707
rect 2053 704 2056 707
rect 2097 704 2102 713
rect 2161 716 2171 720
rect 2216 720 2221 727
rect 2161 712 2165 716
rect 2228 720 2233 727
rect 2313 720 2318 730
rect 2356 727 2404 732
rect 2506 734 2511 740
rect 2543 734 2548 740
rect 2568 741 2684 742
rect 2568 731 2572 741
rect 2633 740 2684 741
rect 2633 734 2638 740
rect 2161 709 2202 712
rect 2161 706 2165 709
rect 2199 706 2202 709
rect 2243 706 2248 715
rect 2308 716 2318 720
rect 2363 720 2368 727
rect 2308 712 2312 716
rect 2375 720 2380 727
rect 2525 719 2530 729
rect 2568 726 2616 731
rect 2642 734 2647 740
rect 2679 734 2684 740
rect 2704 731 2708 742
rect 2779 736 2784 742
rect 2788 736 2793 742
rect 2825 736 2830 742
rect 2850 733 2854 744
rect 2926 742 2977 744
rect 2926 736 2931 742
rect 2308 709 2349 712
rect 1862 683 1909 688
rect 1946 687 1951 691
rect 1998 688 2001 702
rect 2043 699 2045 702
rect 2053 700 2085 704
rect 2097 700 2118 704
rect 2025 696 2028 699
rect 2042 688 2045 699
rect 2097 696 2102 700
rect 1941 682 1976 687
rect 1998 683 2045 688
rect 1872 673 1877 674
rect 1895 673 1900 674
rect 1972 661 1976 682
rect 2082 687 2087 691
rect 2144 690 2147 704
rect 2189 701 2191 704
rect 2199 702 2231 706
rect 2243 702 2264 706
rect 2171 698 2174 701
rect 2188 690 2191 701
rect 2243 698 2248 702
rect 2308 706 2312 709
rect 2346 706 2349 709
rect 2390 706 2395 715
rect 2520 715 2530 719
rect 2575 719 2580 726
rect 2520 711 2524 715
rect 2587 719 2592 726
rect 2661 719 2666 729
rect 2704 726 2752 731
rect 2520 708 2561 711
rect 2077 686 2112 687
rect 2077 682 2125 686
rect 2144 685 2191 690
rect 2228 689 2233 693
rect 2291 690 2294 704
rect 2336 701 2338 704
rect 2346 702 2378 706
rect 2390 702 2420 706
rect 2318 698 2321 701
rect 2335 690 2338 701
rect 2390 698 2395 702
rect 2520 705 2524 708
rect 2558 705 2561 708
rect 2602 705 2607 714
rect 2656 715 2666 719
rect 2711 719 2716 726
rect 2656 711 2660 715
rect 2723 719 2728 726
rect 2807 721 2812 731
rect 2850 728 2898 733
rect 2935 736 2940 742
rect 2972 736 2977 742
rect 2997 733 3001 744
rect 2656 708 2697 711
rect 2656 705 2660 708
rect 2694 705 2697 708
rect 2738 705 2743 714
rect 2802 717 2812 721
rect 2857 721 2862 728
rect 2802 713 2806 717
rect 2869 721 2874 728
rect 2954 721 2959 731
rect 2997 728 3045 733
rect 2802 710 2843 713
rect 2802 707 2806 710
rect 2840 707 2843 710
rect 2884 707 2889 716
rect 2949 717 2959 721
rect 3004 721 3009 728
rect 2949 713 2953 717
rect 3016 721 3021 728
rect 2949 710 2990 713
rect 2949 707 2953 710
rect 2987 707 2990 710
rect 3031 707 3036 716
rect 2223 684 2261 689
rect 2291 685 2338 690
rect 2106 681 2125 682
rect 2008 673 2013 674
rect 2031 673 2036 674
rect 2116 661 2123 681
rect 2154 675 2159 676
rect 2177 675 2182 676
rect 2252 661 2261 684
rect 2375 689 2380 693
rect 2503 689 2506 703
rect 2548 700 2550 703
rect 2558 701 2590 705
rect 2602 701 2610 705
rect 2530 697 2533 700
rect 2547 689 2550 700
rect 2602 697 2607 701
rect 2370 684 2406 689
rect 2503 684 2550 689
rect 2301 675 2306 676
rect 2324 675 2329 676
rect 2397 661 2406 684
rect 2587 688 2592 692
rect 2639 689 2642 703
rect 2684 700 2686 703
rect 2694 701 2726 705
rect 2738 701 2746 705
rect 2666 697 2669 700
rect 2683 689 2686 700
rect 2738 697 2743 701
rect 2582 683 2617 688
rect 2639 684 2686 689
rect 2513 674 2518 675
rect 2536 674 2541 675
rect 2613 662 2617 683
rect 2723 688 2728 692
rect 2785 691 2788 705
rect 2830 702 2832 705
rect 2840 703 2872 707
rect 2884 703 2892 707
rect 2812 699 2815 702
rect 2829 691 2832 702
rect 2884 699 2889 703
rect 2718 687 2753 688
rect 2718 683 2766 687
rect 2785 686 2832 691
rect 2869 690 2874 694
rect 2932 691 2935 705
rect 2977 702 2979 705
rect 2987 703 3019 707
rect 3031 703 3039 707
rect 2959 699 2962 702
rect 2976 691 2979 702
rect 3031 699 3036 703
rect 2864 685 2902 690
rect 2932 686 2979 691
rect 2747 682 2766 683
rect 2649 674 2654 675
rect 2672 674 2677 675
rect 2757 662 2764 682
rect 2795 676 2800 677
rect 2818 676 2823 677
rect 2893 662 2902 685
rect 3016 690 3021 694
rect 3011 685 3047 690
rect 2942 676 2947 677
rect 2965 676 2970 677
rect 3038 662 3047 685
rect 2425 661 2433 662
rect 1972 655 2433 661
rect 2613 657 3048 662
rect 2613 656 3023 657
rect 2425 644 2433 655
rect 2634 644 2643 656
rect 2342 639 2373 640
rect 2197 638 2373 639
rect 1835 636 1865 638
rect 2073 637 2373 638
rect 1904 636 1935 637
rect 2048 636 2373 637
rect 2424 636 2643 644
rect 1835 635 2345 636
rect 1835 633 2200 635
rect 2209 634 2345 635
rect 1835 631 1907 633
rect 1926 631 2051 633
rect 1856 625 1861 631
rect 1865 625 1870 631
rect 1902 625 1907 631
rect 1927 622 1931 631
rect 2000 625 2005 631
rect 1884 610 1889 620
rect 1927 617 1975 622
rect 2009 625 2014 631
rect 2046 625 2051 631
rect 2071 622 2075 633
rect 2149 627 2154 633
rect 2158 627 2163 633
rect 2195 627 2200 633
rect 2220 624 2224 634
rect 2294 628 2299 634
rect 1879 606 1889 610
rect 1934 610 1939 617
rect 1879 602 1883 606
rect 1946 610 1951 617
rect 2028 610 2033 620
rect 2071 617 2119 622
rect 1879 599 1920 602
rect 1879 596 1883 599
rect 1917 596 1920 599
rect 1961 596 1966 605
rect 2023 606 2033 610
rect 2078 610 2083 617
rect 2023 602 2027 606
rect 2090 610 2095 617
rect 2177 612 2182 622
rect 2220 619 2268 624
rect 2303 628 2308 634
rect 2340 628 2345 634
rect 2365 625 2369 636
rect 2023 599 2064 602
rect 1862 580 1865 594
rect 1907 591 1909 594
rect 1917 592 1949 596
rect 1961 592 1993 596
rect 1889 588 1892 591
rect 1906 580 1909 591
rect 1961 588 1966 592
rect 2023 596 2027 599
rect 2061 596 2064 599
rect 2105 596 2110 605
rect 2172 608 2182 612
rect 2227 612 2232 619
rect 2172 604 2176 608
rect 2239 612 2244 619
rect 2322 613 2327 623
rect 2365 620 2413 625
rect 2172 601 2213 604
rect 2172 598 2176 601
rect 2210 598 2213 601
rect 2254 598 2259 607
rect 2317 609 2327 613
rect 2372 613 2377 620
rect 2317 605 2321 609
rect 2384 613 2389 620
rect 2317 602 2358 605
rect 2317 599 2321 602
rect 2355 599 2358 602
rect 2399 599 2404 608
rect 1862 575 1909 580
rect 1946 579 1951 583
rect 2006 580 2009 594
rect 2051 591 2053 594
rect 2061 592 2093 596
rect 2105 592 2133 596
rect 2033 588 2036 591
rect 2050 580 2053 591
rect 2105 588 2110 592
rect 1941 574 1976 579
rect 2006 575 2053 580
rect 1597 566 1700 567
rect 1471 563 1701 566
rect 1471 562 1600 563
rect 1471 522 1476 562
rect 1549 561 1600 562
rect 1549 555 1554 561
rect 1558 555 1563 561
rect 1595 555 1600 561
rect 1620 553 1624 563
rect 1693 553 1701 563
rect 1872 565 1877 566
rect 1895 565 1900 566
rect 1577 540 1582 550
rect 1618 548 1701 553
rect 1572 536 1582 540
rect 1625 541 1630 548
rect 1637 541 1642 548
rect 1572 532 1576 536
rect 1572 529 1613 532
rect 1572 526 1576 529
rect 1610 526 1613 529
rect 1652 527 1657 536
rect 1693 528 1701 548
rect 1617 526 1640 527
rect 716 521 1476 522
rect 720 510 724 521
rect 676 505 724 510
rect 744 519 795 521
rect 744 513 749 519
rect 781 513 786 519
rect 790 513 795 519
rect 867 510 871 521
rect 700 498 705 505
rect 712 498 717 505
rect 762 498 767 508
rect 823 505 871 510
rect 891 519 1476 521
rect 891 513 896 519
rect 928 513 933 519
rect 937 513 942 519
rect 1013 508 1017 519
rect 847 498 852 505
rect 762 494 772 498
rect 685 484 690 493
rect 768 490 772 494
rect 731 487 772 490
rect 731 484 734 487
rect 768 484 772 487
rect 859 498 864 505
rect 909 498 914 508
rect 969 503 1017 508
rect 1037 518 1153 519
rect 1037 517 1088 518
rect 1037 511 1042 517
rect 1074 511 1079 517
rect 1083 511 1088 517
rect 1149 508 1153 518
rect 909 494 919 498
rect 993 496 998 503
rect 667 480 690 484
rect 702 480 734 484
rect 685 476 690 480
rect 742 479 744 482
rect 700 467 705 471
rect 742 468 745 479
rect 759 476 762 479
rect 786 468 789 482
rect 832 484 837 493
rect 915 490 919 494
rect 878 487 919 490
rect 878 484 881 487
rect 915 484 919 487
rect 1005 496 1010 503
rect 1055 496 1060 506
rect 1105 503 1153 508
rect 1173 517 1476 519
rect 1173 511 1178 517
rect 1210 511 1215 517
rect 1218 516 1476 517
rect 1219 511 1224 516
rect 1129 496 1134 503
rect 1055 492 1065 496
rect 821 481 837 484
rect 819 480 837 481
rect 849 480 881 484
rect 832 476 837 480
rect 889 479 891 482
rect 674 465 710 467
rect 523 462 710 465
rect 523 460 683 462
rect 742 463 789 468
rect 847 467 852 471
rect 889 468 892 479
rect 906 476 909 479
rect 933 468 936 482
rect 978 482 983 491
rect 1061 488 1065 492
rect 1024 485 1065 488
rect 1024 482 1027 485
rect 1061 482 1065 485
rect 1141 496 1146 503
rect 1191 496 1196 506
rect 1191 492 1201 496
rect 1114 482 1119 491
rect 1197 488 1201 492
rect 1160 485 1201 488
rect 1160 482 1163 485
rect 1197 482 1201 485
rect 966 478 983 482
rect 995 478 1027 482
rect 978 474 983 478
rect 1035 477 1037 480
rect 1104 481 1119 482
rect 819 462 857 467
rect 489 439 494 443
rect 280 430 448 431
rect 474 430 479 434
rect 523 430 529 460
rect 280 426 529 430
rect 443 425 529 426
rect 235 417 404 422
rect 399 412 404 417
rect 421 412 426 416
rect 160 401 198 405
rect 399 407 426 412
rect 160 400 202 401
rect 483 348 488 360
rect 144 343 149 348
rect 379 343 516 348
rect 1 339 149 343
rect 153 339 372 343
rect 1 338 49 339
rect 25 331 30 338
rect 37 331 42 338
rect 57 327 62 339
rect 10 317 15 326
rect 69 327 74 339
rect 101 327 106 339
rect 133 327 138 339
rect 85 319 90 322
rect 70 318 90 319
rect 117 318 122 322
rect 3 313 15 317
rect 27 313 46 317
rect 10 309 15 313
rect 25 300 30 304
rect 42 305 46 313
rect 70 314 122 318
rect 70 305 75 314
rect 42 300 45 305
rect 50 300 75 305
rect 153 305 158 339
rect 168 327 356 331
rect 168 326 308 327
rect 168 319 173 326
rect 205 319 210 326
rect 279 319 284 326
rect 220 305 225 314
rect 291 319 296 326
rect 303 315 308 326
rect 264 305 269 314
rect 315 315 320 327
rect 153 302 208 305
rect 204 301 208 302
rect 220 301 228 305
rect 0 295 39 300
rect 34 279 39 295
rect 70 293 75 300
rect 220 297 225 301
rect 238 301 269 305
rect 281 303 302 305
rect 281 301 288 303
rect 205 288 210 292
rect 133 286 138 288
rect 171 286 227 288
rect 133 283 227 286
rect 133 282 175 283
rect 133 279 138 282
rect 34 275 138 279
rect 153 268 186 271
rect 109 249 114 265
rect 125 260 130 265
rect 125 256 226 260
rect 109 245 143 249
rect 238 237 242 301
rect 264 297 269 301
rect 293 301 302 303
rect 298 298 302 301
rect 349 304 354 310
rect 367 304 372 339
rect 379 341 384 343
rect 398 321 451 327
rect 398 315 403 321
rect 432 304 437 310
rect 349 299 437 304
rect 298 293 319 298
rect 279 288 284 292
rect 255 283 293 288
rect 283 246 288 283
rect 349 276 354 299
rect 398 293 401 296
rect 304 265 309 268
rect 391 288 406 293
rect 383 275 388 288
rect 315 246 320 271
rect 398 276 403 288
rect 432 276 437 299
rect 446 246 451 321
rect 463 283 506 288
rect 465 276 470 283
rect 477 276 482 283
rect 492 263 497 271
rect 511 263 516 343
rect 477 258 480 262
rect 492 258 516 263
rect 492 254 497 258
rect 283 245 451 246
rect 477 245 482 249
rect 523 245 529 425
rect 541 432 542 441
rect 647 439 655 440
rect 674 439 683 460
rect 751 453 756 454
rect 774 453 779 454
rect 819 439 828 462
rect 889 463 936 468
rect 993 465 998 469
rect 1035 466 1038 477
rect 1052 474 1055 477
rect 1079 466 1082 480
rect 1109 478 1119 481
rect 1131 478 1163 482
rect 1114 474 1119 478
rect 1171 477 1173 480
rect 968 464 1003 465
rect 955 460 1003 464
rect 898 453 903 454
rect 955 459 974 460
rect 1035 461 1082 466
rect 1129 465 1134 469
rect 1171 466 1174 477
rect 1188 474 1191 477
rect 1215 466 1218 480
rect 1104 460 1139 465
rect 921 453 926 454
rect 957 439 964 459
rect 1044 451 1049 452
rect 1067 451 1072 452
rect 1104 439 1108 460
rect 1171 461 1218 466
rect 1180 451 1185 452
rect 1203 451 1208 452
rect 541 389 548 432
rect 575 355 581 438
rect 647 433 1108 439
rect 545 349 581 355
rect 618 324 620 333
rect 618 256 627 324
rect 283 241 531 245
rect 446 240 531 241
rect 238 232 407 237
rect 402 227 407 232
rect 424 227 429 231
rect 402 222 429 227
rect 502 203 506 225
rect 379 168 510 173
rect 178 164 372 168
rect 178 130 183 164
rect 193 152 356 156
rect 193 151 308 152
rect 193 144 198 151
rect 205 144 210 151
rect 279 144 284 151
rect 220 130 225 139
rect 291 144 296 151
rect 303 140 308 151
rect 264 130 269 139
rect 315 140 320 152
rect 178 127 208 130
rect 204 126 208 127
rect 220 126 228 130
rect 220 122 225 126
rect 238 126 269 130
rect 281 128 302 130
rect 281 126 288 128
rect 205 113 210 117
rect 196 108 227 113
rect 238 62 242 126
rect 264 122 269 126
rect 294 126 302 128
rect 298 123 302 126
rect 349 129 354 135
rect 367 129 372 164
rect 379 166 384 168
rect 398 146 451 152
rect 398 140 403 146
rect 432 129 437 135
rect 349 124 437 129
rect 298 118 319 123
rect 279 113 284 117
rect 255 108 293 113
rect 283 71 288 108
rect 349 101 354 124
rect 398 118 401 121
rect 388 113 406 118
rect 304 90 309 93
rect 379 101 386 113
rect 398 101 403 113
rect 379 96 383 101
rect 432 101 437 124
rect 315 71 320 96
rect 446 71 451 146
rect 463 108 506 113
rect 465 101 470 108
rect 477 101 482 108
rect 492 88 497 96
rect 511 88 516 168
rect 477 83 480 87
rect 492 83 516 88
rect 492 79 497 83
rect 283 70 451 71
rect 477 70 482 74
rect 523 70 529 240
rect 617 172 627 256
rect 617 107 626 172
rect 283 66 529 70
rect 446 65 529 66
rect 238 57 407 62
rect 402 52 407 57
rect 424 52 429 56
rect 402 47 429 52
rect 476 29 483 38
rect 635 29 641 373
rect 647 327 655 433
rect 707 417 738 418
rect 707 416 883 417
rect 1237 416 1245 516
rect 707 415 1007 416
rect 707 414 1032 415
rect 1145 414 1176 415
rect 1215 414 1245 416
rect 1471 414 1476 516
rect 1555 510 1558 524
rect 1600 521 1602 524
rect 1610 523 1640 526
rect 1652 523 1660 527
rect 1610 522 1637 523
rect 1582 518 1585 521
rect 1599 510 1602 521
rect 1652 519 1657 523
rect 1694 523 1700 528
rect 1834 523 1837 553
rect 1968 550 1977 574
rect 2090 579 2095 583
rect 2155 582 2158 596
rect 2200 593 2202 596
rect 2210 594 2242 598
rect 2254 594 2282 598
rect 2182 590 2185 593
rect 2199 582 2202 593
rect 2254 590 2259 594
rect 2085 574 2126 579
rect 2155 577 2202 582
rect 2239 581 2244 585
rect 2300 583 2303 597
rect 2345 594 2347 597
rect 2355 595 2387 599
rect 2399 595 2407 599
rect 2327 591 2330 594
rect 2344 583 2347 594
rect 2399 591 2404 595
rect 2234 576 2269 581
rect 2300 578 2347 583
rect 2384 582 2389 586
rect 2408 582 2415 583
rect 2379 577 2415 582
rect 2016 565 2021 566
rect 2039 565 2044 566
rect 2118 550 2125 574
rect 2165 567 2170 568
rect 2188 567 2193 568
rect 2262 550 2269 576
rect 2310 567 2315 569
rect 2333 568 2338 569
rect 2408 550 2415 577
rect 1968 549 2415 550
rect 2425 549 2433 636
rect 2634 635 2643 636
rect 1968 544 2433 549
rect 1637 510 1642 514
rect 1555 505 1602 510
rect 1634 505 1656 510
rect 1649 504 1656 505
rect 711 403 715 414
rect 667 398 715 403
rect 735 413 1245 414
rect 735 412 871 413
rect 735 406 740 412
rect 772 406 777 412
rect 781 406 786 412
rect 856 402 860 412
rect 691 391 696 398
rect 703 391 708 398
rect 753 391 758 401
rect 812 397 860 402
rect 880 411 1245 413
rect 880 405 885 411
rect 917 405 922 411
rect 926 405 931 411
rect 1005 400 1009 411
rect 753 387 763 391
rect 836 390 841 397
rect 676 377 681 386
rect 759 383 763 387
rect 722 380 763 383
rect 722 377 725 380
rect 759 377 763 380
rect 848 390 853 397
rect 898 390 903 400
rect 961 395 1009 400
rect 1029 409 1154 411
rect 1173 409 1245 411
rect 1390 409 1476 414
rect 1693 509 1701 523
rect 1692 504 1702 509
rect 1029 403 1034 409
rect 1066 403 1071 409
rect 1075 403 1080 409
rect 1149 400 1153 409
rect 898 386 908 390
rect 985 388 990 395
rect 668 373 681 377
rect 693 373 725 377
rect 676 369 681 373
rect 733 372 735 375
rect 665 360 672 361
rect 691 360 696 364
rect 733 361 736 372
rect 750 369 753 372
rect 777 361 780 375
rect 821 376 826 385
rect 904 382 908 386
rect 867 379 908 382
rect 867 376 870 379
rect 904 376 908 379
rect 997 388 1002 395
rect 1047 388 1052 398
rect 1105 395 1153 400
rect 1173 403 1178 409
rect 1210 403 1215 409
rect 1219 403 1224 409
rect 1397 402 1402 409
rect 1129 388 1134 395
rect 1047 384 1057 388
rect 809 373 826 376
rect 818 372 826 373
rect 838 372 870 376
rect 821 368 826 372
rect 878 371 880 374
rect 970 374 975 383
rect 1053 380 1057 384
rect 1016 377 1057 380
rect 1016 374 1019 377
rect 1053 374 1057 377
rect 1141 388 1146 395
rect 1191 388 1196 398
rect 1409 402 1414 409
rect 1447 402 1452 409
rect 1191 384 1201 388
rect 665 355 701 360
rect 665 328 672 355
rect 733 356 780 361
rect 836 359 841 363
rect 878 360 881 371
rect 895 368 898 371
rect 922 360 925 374
rect 952 369 975 374
rect 987 370 1019 374
rect 970 366 975 369
rect 1027 369 1029 372
rect 811 354 846 359
rect 742 346 747 347
rect 765 345 770 347
rect 811 328 818 354
rect 878 355 925 360
rect 985 357 990 361
rect 1027 358 1030 369
rect 1044 366 1047 369
rect 1071 358 1074 372
rect 1114 374 1119 383
rect 1197 380 1201 384
rect 1410 384 1412 388
rect 1410 383 1411 384
rect 1424 380 1429 397
rect 1462 388 1467 397
rect 1447 384 1450 388
rect 1462 383 1465 388
rect 1462 380 1467 383
rect 1160 377 1201 380
rect 1160 374 1163 377
rect 1197 374 1201 377
rect 1095 370 1119 374
rect 1131 370 1163 374
rect 1114 366 1119 370
rect 1171 369 1173 372
rect 954 352 995 357
rect 887 345 892 346
rect 910 345 915 346
rect 955 328 962 352
rect 1027 353 1074 358
rect 1129 357 1134 361
rect 1171 358 1174 369
rect 1188 366 1191 369
rect 1215 358 1218 372
rect 1409 371 1414 375
rect 1447 373 1452 375
rect 1434 371 1453 373
rect 1353 370 1479 371
rect 1353 366 1437 370
rect 1450 368 1479 370
rect 1452 366 1479 368
rect 1353 363 1404 366
rect 1104 352 1139 357
rect 1036 343 1041 344
rect 1059 343 1064 344
rect 1103 328 1112 352
rect 1171 353 1218 358
rect 1180 343 1185 344
rect 1203 343 1208 344
rect 1249 335 1318 339
rect 665 327 1112 328
rect 647 322 1112 327
rect 665 321 672 322
rect 955 320 962 322
rect 1103 303 1111 322
rect 1398 303 1404 363
rect 1103 299 1405 303
rect 1319 131 1323 171
rect 1398 161 1404 299
rect 1442 262 1446 361
rect 1488 274 1496 482
rect 1596 448 1627 449
rect 1548 445 1627 448
rect 1548 443 1599 445
rect 1548 437 1553 443
rect 1557 437 1562 443
rect 1594 437 1599 443
rect 1619 434 1623 445
rect 1693 434 1701 504
rect 1935 509 1944 511
rect 1729 504 1944 509
rect 1576 422 1581 432
rect 1617 429 1701 434
rect 1571 418 1581 422
rect 1624 422 1629 429
rect 1571 414 1575 418
rect 1636 422 1641 429
rect 1674 428 1688 429
rect 1571 411 1612 414
rect 1571 408 1575 411
rect 1609 408 1612 411
rect 1651 408 1656 417
rect 1554 392 1557 406
rect 1599 403 1601 406
rect 1609 404 1639 408
rect 1651 404 1666 408
rect 1581 400 1584 403
rect 1598 392 1601 403
rect 1651 400 1656 404
rect 1554 387 1601 392
rect 1636 391 1641 395
rect 1632 386 1662 391
rect 1564 375 1569 378
rect 1586 375 1592 378
rect 1693 380 1701 429
rect 1792 427 1796 485
rect 1855 476 1891 481
rect 1888 460 1891 476
rect 1935 475 1944 504
rect 2076 475 2083 544
rect 2118 542 2125 544
rect 2408 543 2415 544
rect 1935 469 2084 475
rect 2076 467 2083 469
rect 2162 465 2388 467
rect 2162 464 2383 465
rect 2162 460 2165 464
rect 1888 457 2165 460
rect 2587 458 2687 459
rect 2734 458 2765 459
rect 2539 457 2765 458
rect 2305 456 2336 457
rect 2441 456 2765 457
rect 2236 455 2765 456
rect 2236 453 2590 455
rect 2236 451 2308 453
rect 2236 450 2263 451
rect 1792 424 2222 427
rect 1738 408 2032 409
rect 1738 407 2042 408
rect 1738 404 2036 407
rect 2024 401 2036 404
rect 2218 399 2222 424
rect 2236 381 2244 450
rect 2257 445 2262 450
rect 2266 445 2271 451
rect 2303 445 2308 451
rect 2328 452 2444 453
rect 2328 442 2332 452
rect 2393 451 2444 452
rect 2393 445 2398 451
rect 2285 430 2290 440
rect 2328 437 2376 442
rect 2402 445 2407 451
rect 2439 445 2444 451
rect 2464 442 2468 453
rect 2539 447 2544 453
rect 2548 447 2553 453
rect 2585 447 2590 453
rect 2610 444 2614 455
rect 2686 453 2737 455
rect 2686 447 2691 453
rect 2280 426 2290 430
rect 2335 430 2340 437
rect 2280 422 2284 426
rect 2347 430 2352 437
rect 2421 430 2426 440
rect 2464 437 2512 442
rect 2280 419 2321 422
rect 2280 416 2284 419
rect 2318 416 2321 419
rect 2362 416 2367 425
rect 2416 426 2426 430
rect 2471 430 2476 437
rect 2416 422 2420 426
rect 2483 430 2488 437
rect 2567 432 2572 442
rect 2610 439 2658 444
rect 2695 447 2700 453
rect 2732 447 2737 453
rect 2757 444 2761 455
rect 2416 419 2457 422
rect 2416 416 2420 419
rect 2454 416 2457 419
rect 2498 416 2503 425
rect 2562 428 2572 432
rect 2617 432 2622 439
rect 2562 424 2566 428
rect 2629 432 2634 439
rect 2714 432 2719 442
rect 2757 439 2805 444
rect 2562 421 2603 424
rect 2562 418 2566 421
rect 2600 418 2603 421
rect 2644 418 2649 427
rect 2709 428 2719 432
rect 2764 432 2769 439
rect 2709 424 2713 428
rect 2776 432 2781 439
rect 2709 421 2750 424
rect 2709 418 2713 421
rect 2747 418 2750 421
rect 2791 418 2796 427
rect 2263 400 2266 414
rect 2308 411 2310 414
rect 2318 412 2350 416
rect 2362 412 2370 416
rect 2290 408 2293 411
rect 2307 400 2310 411
rect 2362 408 2367 412
rect 2263 395 2310 400
rect 2347 399 2352 403
rect 2399 400 2402 414
rect 2444 411 2446 414
rect 2454 412 2486 416
rect 2498 412 2506 416
rect 2426 408 2429 411
rect 2443 400 2446 411
rect 2498 408 2503 412
rect 2342 394 2377 399
rect 2399 395 2446 400
rect 2055 380 2244 381
rect 1693 376 2244 380
rect 2273 385 2278 386
rect 2296 385 2301 386
rect 1693 375 2055 376
rect 1595 344 1626 345
rect 1547 341 1626 344
rect 1547 339 1598 341
rect 1547 333 1552 339
rect 1556 333 1561 339
rect 1593 333 1598 339
rect 1618 330 1622 341
rect 1693 330 1701 375
rect 1995 367 2000 375
rect 1769 362 1984 366
rect 2005 367 2010 375
rect 2062 369 2067 376
rect 2024 362 2029 367
rect 2074 369 2079 376
rect 1980 352 1984 362
rect 1980 348 2008 352
rect 2004 347 2008 348
rect 2043 351 2048 362
rect 2089 355 2094 364
rect 2061 351 2077 355
rect 2089 351 2099 355
rect 2043 346 2065 351
rect 2089 347 2094 351
rect 2043 344 2048 346
rect 1575 318 1580 328
rect 1618 325 1701 330
rect 2005 338 2048 344
rect 2236 350 2244 376
rect 2373 373 2377 394
rect 2483 399 2488 403
rect 2545 402 2548 416
rect 2590 413 2592 416
rect 2600 414 2632 418
rect 2644 414 2652 418
rect 2572 410 2575 413
rect 2589 402 2592 413
rect 2644 410 2649 414
rect 2478 398 2513 399
rect 2478 394 2526 398
rect 2545 397 2592 402
rect 2629 401 2634 405
rect 2692 402 2695 416
rect 2737 413 2739 416
rect 2747 414 2779 418
rect 2791 414 2799 418
rect 2719 410 2722 413
rect 2736 402 2739 413
rect 2791 410 2796 414
rect 2624 396 2662 401
rect 2692 397 2739 402
rect 2507 393 2526 394
rect 2409 385 2414 386
rect 2432 385 2437 386
rect 2517 373 2524 393
rect 2555 387 2560 388
rect 2578 387 2583 388
rect 2653 373 2662 396
rect 2776 401 2781 405
rect 2771 396 2807 401
rect 2702 387 2707 388
rect 2725 387 2730 388
rect 2798 373 2807 396
rect 2826 373 2834 374
rect 2373 367 2834 373
rect 2743 351 2774 352
rect 2598 350 2774 351
rect 2236 348 2266 350
rect 2474 349 2774 350
rect 2305 348 2336 349
rect 2449 348 2774 349
rect 2236 347 2746 348
rect 2236 345 2601 347
rect 2610 346 2746 347
rect 2236 343 2308 345
rect 2327 343 2452 345
rect 2074 338 2079 342
rect 2005 330 2010 338
rect 2043 330 2048 338
rect 2065 337 2104 338
rect 2257 337 2262 343
rect 2065 333 2243 337
rect 1570 314 1580 318
rect 1625 318 1630 325
rect 1570 310 1574 314
rect 1637 318 1642 325
rect 1570 307 1611 310
rect 1570 304 1574 307
rect 1608 304 1611 307
rect 1652 304 1657 313
rect 1553 288 1556 302
rect 1598 299 1600 302
rect 1608 300 1640 304
rect 1652 300 1670 304
rect 1580 296 1583 299
rect 1597 288 1600 299
rect 1652 296 1657 300
rect 1553 283 1600 288
rect 1637 287 1642 291
rect 1631 282 1658 287
rect 1488 269 1568 274
rect 1586 262 1591 274
rect 1442 256 1591 262
rect 1533 179 1537 256
rect 1595 248 1626 249
rect 1547 245 1626 248
rect 1547 243 1598 245
rect 1547 237 1552 243
rect 1556 237 1561 243
rect 1593 237 1598 243
rect 1618 234 1622 245
rect 1693 234 1701 325
rect 2023 319 2028 325
rect 2065 319 2070 333
rect 2100 332 2243 333
rect 2266 337 2271 343
rect 2303 337 2308 343
rect 2328 334 2332 343
rect 2401 337 2406 343
rect 2023 316 2070 319
rect 2028 312 2032 316
rect 1616 233 1701 234
rect 2019 309 2032 312
rect 1575 222 1580 232
rect 1616 229 2002 233
rect 1570 218 1580 222
rect 1624 222 1629 229
rect 1570 214 1574 218
rect 1636 222 1641 229
rect 1687 228 2002 229
rect 1570 211 1611 214
rect 1570 208 1574 211
rect 1608 208 1611 211
rect 1651 208 1656 217
rect 1553 192 1556 206
rect 1598 203 1600 206
rect 1608 204 1639 208
rect 1651 204 1805 208
rect 1580 200 1583 203
rect 1597 192 1600 203
rect 1651 200 1656 204
rect 1553 187 1600 192
rect 1636 191 1641 195
rect 1657 191 1665 192
rect 1632 186 1665 191
rect 1657 185 1665 186
rect 1774 185 1938 188
rect 1533 178 1563 179
rect 1533 175 1568 178
rect 1659 161 1665 185
rect 1398 160 1665 161
rect 1398 156 2006 160
rect 2019 160 2023 309
rect 2238 254 2243 332
rect 2285 322 2290 332
rect 2328 329 2376 334
rect 2410 337 2415 343
rect 2447 337 2452 343
rect 2472 334 2476 345
rect 2550 339 2555 345
rect 2559 339 2564 345
rect 2596 339 2601 345
rect 2621 336 2625 346
rect 2695 340 2700 346
rect 2280 318 2290 322
rect 2335 322 2340 329
rect 2280 314 2284 318
rect 2347 322 2352 329
rect 2429 322 2434 332
rect 2472 329 2520 334
rect 2280 311 2321 314
rect 2280 308 2284 311
rect 2318 308 2321 311
rect 2263 292 2266 306
rect 2308 303 2310 306
rect 2318 304 2350 308
rect 2290 300 2293 303
rect 2307 292 2310 303
rect 2362 300 2367 317
rect 2424 318 2434 322
rect 2479 322 2484 329
rect 2424 314 2428 318
rect 2491 322 2496 329
rect 2578 324 2583 334
rect 2621 331 2669 336
rect 2704 340 2709 346
rect 2741 340 2746 346
rect 2766 337 2770 348
rect 2424 311 2465 314
rect 2424 308 2428 311
rect 2462 308 2465 311
rect 2506 308 2511 317
rect 2573 320 2583 324
rect 2628 324 2633 331
rect 2573 316 2577 320
rect 2640 324 2645 331
rect 2723 325 2728 335
rect 2766 332 2814 337
rect 2573 313 2614 316
rect 2573 310 2577 313
rect 2611 310 2614 313
rect 2655 310 2660 319
rect 2718 321 2728 325
rect 2773 325 2778 332
rect 2718 317 2722 321
rect 2785 325 2790 332
rect 2718 314 2759 317
rect 2718 311 2722 314
rect 2756 311 2759 314
rect 2800 311 2805 320
rect 2263 287 2310 292
rect 2347 291 2352 295
rect 2407 292 2410 306
rect 2452 303 2454 306
rect 2462 304 2494 308
rect 2506 304 2520 308
rect 2434 300 2437 303
rect 2451 292 2454 303
rect 2506 300 2511 304
rect 2342 286 2377 291
rect 2407 287 2454 292
rect 2273 277 2278 278
rect 2296 277 2301 278
rect 2369 262 2378 286
rect 2491 291 2496 295
rect 2556 294 2559 308
rect 2601 305 2603 308
rect 2611 306 2643 310
rect 2655 306 2667 310
rect 2583 302 2586 305
rect 2600 294 2603 305
rect 2655 302 2660 306
rect 2486 286 2527 291
rect 2556 289 2603 294
rect 2640 293 2645 297
rect 2701 295 2704 309
rect 2746 306 2748 309
rect 2756 307 2788 311
rect 2800 307 2812 311
rect 2728 303 2731 306
rect 2745 295 2748 306
rect 2800 303 2805 307
rect 2635 288 2670 293
rect 2701 290 2748 295
rect 2785 294 2790 298
rect 2809 294 2816 295
rect 2780 289 2816 294
rect 2417 277 2422 278
rect 2440 277 2445 278
rect 2519 262 2526 286
rect 2566 279 2571 280
rect 2589 279 2594 280
rect 2663 262 2670 288
rect 2711 279 2716 281
rect 2734 280 2739 281
rect 2809 262 2816 289
rect 2369 261 2816 262
rect 2826 261 2834 367
rect 2369 256 2834 261
rect 2369 254 2375 256
rect 2519 254 2526 256
rect 2809 255 2816 256
rect 2238 251 2375 254
rect 2011 156 2023 160
rect 2135 138 2272 143
rect 2135 136 2140 138
rect 1319 126 1831 131
rect 2007 122 2036 126
rect 2042 122 2112 126
rect 2007 121 2055 122
rect 2031 114 2036 121
rect 2043 114 2048 121
rect 2059 110 2064 122
rect 2016 100 2021 109
rect 2071 110 2076 122
rect 2154 116 2207 122
rect 2154 110 2159 116
rect 1994 96 2021 100
rect 2033 96 2046 100
rect 476 23 641 29
rect 673 6 682 92
rect 1994 32 1998 96
rect 2016 92 2021 96
rect 2051 96 2058 100
rect 2054 93 2058 96
rect 2105 99 2110 105
rect 2188 99 2193 105
rect 2105 94 2193 99
rect 2054 88 2075 93
rect 2031 83 2036 87
rect 2012 78 2045 83
rect 2039 41 2044 78
rect 2105 71 2110 94
rect 2154 88 2157 91
rect 2152 83 2162 88
rect 2060 60 2065 63
rect 2154 71 2159 83
rect 2071 41 2076 66
rect 2188 71 2193 94
rect 2202 41 2207 116
rect 2219 78 2262 83
rect 2221 71 2226 78
rect 2233 71 2238 78
rect 2248 58 2253 66
rect 2267 58 2272 138
rect 2233 53 2236 57
rect 2248 53 2272 58
rect 2248 49 2253 53
rect 2039 40 2207 41
rect 2233 40 2238 44
rect 2039 36 2263 40
rect 2202 35 2263 36
rect 1994 27 2163 32
rect 2158 22 2163 27
rect 2180 22 2185 26
rect 1459 15 1601 20
rect 2158 17 2185 22
rect 1483 8 1488 15
rect 299 0 682 6
rect 1495 8 1500 15
rect 1522 4 1527 15
rect 1579 4 1584 15
rect 1468 -6 1473 3
rect 1422 -10 1473 -6
rect 1485 -10 1511 -6
rect 1468 -14 1473 -10
rect 1483 -23 1488 -19
rect 1508 -23 1511 -10
rect 1531 -23 1536 -1
rect 1458 -28 1505 -23
rect 1508 -27 1568 -23
rect 1500 -40 1505 -28
rect 1531 -32 1536 -27
rect 1563 -32 1568 -27
rect 1547 -40 1552 -37
rect 1500 -41 1552 -40
rect 1579 -40 1584 -37
rect 1500 -44 1579 -41
rect 1539 -56 1544 -55
rect 1555 -57 1560 -55
rect 1571 -57 1576 -55
rect 1328 -99 1356 -98
rect 1328 -100 1404 -99
rect 1328 -101 1502 -100
rect 1595 -101 1601 15
rect 2129 -45 2266 -40
rect 2129 -47 2134 -45
rect 2001 -61 2106 -57
rect 2001 -62 2049 -61
rect 2025 -69 2030 -62
rect 2053 -73 2058 -61
rect 2010 -83 2015 -74
rect 2065 -73 2070 -61
rect 2148 -67 2201 -61
rect 2148 -73 2153 -67
rect 1988 -87 2015 -83
rect 2027 -87 2038 -83
rect 2043 -87 2052 -83
rect 1607 -101 1638 -100
rect 1834 -101 1839 -100
rect 1328 -102 1839 -101
rect 1329 -113 1333 -102
rect 1259 -117 1333 -113
rect 1353 -104 1839 -102
rect 1353 -110 1358 -104
rect 1390 -110 1395 -104
rect 1399 -110 1404 -104
rect 1475 -115 1479 -104
rect 1234 -202 1239 -148
rect 1259 -217 1265 -117
rect 1285 -118 1333 -117
rect 1309 -125 1314 -118
rect 1321 -125 1326 -118
rect 1371 -125 1376 -115
rect 1431 -120 1479 -115
rect 1499 -105 1615 -104
rect 1499 -106 1550 -105
rect 1499 -112 1504 -106
rect 1536 -112 1541 -106
rect 1545 -112 1550 -106
rect 1611 -115 1615 -105
rect 1371 -129 1381 -125
rect 1455 -127 1460 -120
rect 1294 -139 1299 -130
rect 1377 -133 1381 -129
rect 1340 -136 1381 -133
rect 1340 -139 1343 -136
rect 1377 -139 1381 -136
rect 1467 -127 1472 -120
rect 1517 -127 1522 -117
rect 1567 -120 1615 -115
rect 1635 -106 1839 -104
rect 1635 -112 1640 -106
rect 1672 -112 1677 -106
rect 1680 -107 1839 -106
rect 1681 -112 1686 -107
rect 1591 -127 1596 -120
rect 1517 -131 1527 -127
rect 1276 -143 1299 -139
rect 1311 -143 1343 -139
rect 1294 -147 1299 -143
rect 1351 -144 1353 -141
rect 1309 -156 1314 -152
rect 1351 -155 1354 -144
rect 1368 -147 1371 -144
rect 1395 -155 1398 -141
rect 1440 -141 1445 -132
rect 1523 -135 1527 -131
rect 1486 -138 1527 -135
rect 1486 -141 1489 -138
rect 1523 -141 1527 -138
rect 1603 -127 1608 -120
rect 1653 -127 1658 -117
rect 1653 -131 1663 -127
rect 1423 -145 1445 -141
rect 1457 -145 1489 -141
rect 1440 -149 1445 -145
rect 1497 -146 1499 -143
rect 1281 -161 1319 -156
rect 1281 -181 1290 -161
rect 1351 -160 1398 -155
rect 1455 -158 1460 -154
rect 1497 -157 1500 -146
rect 1514 -149 1517 -146
rect 1541 -157 1544 -143
rect 1576 -141 1581 -132
rect 1659 -135 1663 -131
rect 1622 -138 1663 -135
rect 1622 -141 1625 -138
rect 1659 -141 1663 -138
rect 1564 -145 1581 -141
rect 1593 -145 1625 -141
rect 1576 -149 1581 -145
rect 1633 -146 1635 -143
rect 1430 -159 1465 -158
rect 1417 -163 1465 -159
rect 1360 -170 1365 -169
rect 1417 -164 1436 -163
rect 1497 -162 1544 -157
rect 1591 -158 1596 -154
rect 1633 -157 1636 -146
rect 1650 -149 1653 -146
rect 1677 -157 1680 -143
rect 1566 -163 1601 -158
rect 1383 -170 1388 -169
rect 1419 -184 1426 -164
rect 1506 -172 1511 -171
rect 1529 -172 1534 -171
rect 1566 -184 1570 -163
rect 1633 -162 1680 -157
rect 1642 -172 1647 -171
rect 1665 -172 1670 -171
rect 1290 -188 1570 -184
rect 1280 -189 1570 -188
rect 1289 -208 1290 -203
rect 1441 -208 1446 -198
rect 1700 -193 1785 -192
rect 1647 -196 1785 -193
rect 1647 -197 1704 -196
rect 1642 -208 1647 -198
rect 1282 -214 1446 -208
rect 1223 -234 1360 -229
rect 1441 -230 1446 -214
rect 1223 -314 1228 -234
rect 1355 -236 1360 -234
rect 1552 -213 1647 -208
rect 1288 -256 1341 -250
rect 1383 -250 1500 -246
rect 1233 -294 1276 -289
rect 1257 -301 1262 -294
rect 1269 -301 1274 -294
rect 1242 -314 1247 -306
rect 1223 -319 1247 -314
rect 1259 -319 1262 -315
rect 1242 -323 1247 -319
rect 1257 -332 1262 -328
rect 1288 -331 1293 -256
rect 1336 -262 1341 -256
rect 1419 -262 1424 -250
rect 1431 -262 1436 -250
rect 1451 -251 1500 -250
rect 1455 -258 1460 -251
rect 1467 -258 1472 -251
rect 1302 -273 1307 -267
rect 1302 -278 1366 -273
rect 1385 -273 1390 -267
rect 1482 -272 1487 -263
rect 1372 -278 1390 -273
rect 1302 -301 1307 -278
rect 1338 -284 1341 -281
rect 1333 -289 1343 -284
rect 1336 -301 1341 -289
rect 1385 -301 1390 -278
rect 1437 -279 1441 -272
rect 1446 -276 1470 -272
rect 1482 -276 1501 -272
rect 1420 -284 1441 -279
rect 1482 -280 1487 -276
rect 1467 -289 1472 -285
rect 1451 -294 1492 -289
rect 1419 -331 1424 -306
rect 1430 -312 1435 -309
rect 1451 -331 1456 -294
rect 1288 -332 1451 -331
rect 1236 -336 1451 -332
rect 1236 -337 1293 -336
rect 1497 -340 1501 -276
rect 1310 -350 1315 -346
rect 1332 -345 1501 -340
rect 1552 -344 1557 -213
rect 1561 -234 1698 -229
rect 1561 -314 1566 -234
rect 1693 -236 1698 -234
rect 1834 -246 1839 -107
rect 1988 -151 1992 -87
rect 2010 -91 2015 -87
rect 2048 -90 2052 -87
rect 2099 -84 2104 -78
rect 2182 -84 2187 -78
rect 2099 -89 2187 -84
rect 2048 -95 2069 -90
rect 2025 -100 2030 -96
rect 2004 -105 2039 -100
rect 2033 -142 2038 -105
rect 2099 -112 2104 -89
rect 2148 -95 2151 -92
rect 2146 -100 2156 -95
rect 2054 -123 2059 -120
rect 2148 -112 2153 -100
rect 2065 -142 2070 -117
rect 2182 -112 2187 -89
rect 2196 -142 2201 -67
rect 2213 -105 2256 -100
rect 2215 -112 2220 -105
rect 2227 -112 2232 -105
rect 2242 -125 2247 -117
rect 2261 -125 2266 -45
rect 2227 -130 2230 -126
rect 2242 -130 2266 -125
rect 2242 -134 2247 -130
rect 2033 -143 2201 -142
rect 2227 -143 2232 -139
rect 2033 -147 2257 -143
rect 2196 -148 2257 -147
rect 1988 -156 2157 -151
rect 2152 -161 2157 -156
rect 2174 -161 2179 -157
rect 2152 -166 2179 -161
rect 2117 -217 2254 -212
rect 2117 -219 2122 -217
rect 1989 -233 2094 -229
rect 1989 -234 2037 -233
rect 2013 -241 2018 -234
rect 1626 -256 1679 -250
rect 1721 -250 1839 -246
rect 1571 -294 1614 -289
rect 1595 -301 1600 -294
rect 1607 -301 1612 -294
rect 1580 -314 1585 -306
rect 1561 -319 1585 -314
rect 1597 -319 1600 -315
rect 1580 -323 1585 -319
rect 1595 -332 1600 -328
rect 1626 -331 1631 -256
rect 1674 -262 1679 -256
rect 1757 -262 1762 -250
rect 1769 -262 1774 -250
rect 1784 -251 1839 -250
rect 2041 -245 2046 -233
rect 1787 -258 1792 -251
rect 1799 -258 1804 -251
rect 1998 -255 2003 -246
rect 2053 -245 2058 -233
rect 2136 -239 2189 -233
rect 2136 -245 2141 -239
rect 1640 -273 1645 -267
rect 1723 -273 1728 -267
rect 1814 -272 1819 -263
rect 1976 -259 2003 -255
rect 2015 -259 2027 -255
rect 2032 -259 2040 -255
rect 1640 -278 1706 -273
rect 1711 -278 1728 -273
rect 1640 -301 1645 -278
rect 1676 -284 1679 -281
rect 1671 -289 1681 -284
rect 1674 -301 1679 -289
rect 1723 -301 1728 -278
rect 1775 -279 1779 -272
rect 1784 -276 1802 -272
rect 1814 -276 1839 -272
rect 1758 -284 1779 -279
rect 1814 -280 1819 -276
rect 1799 -289 1804 -285
rect 1789 -294 1829 -289
rect 1757 -331 1762 -306
rect 1768 -312 1773 -309
rect 1789 -331 1794 -294
rect 1626 -332 1794 -331
rect 1577 -336 1794 -332
rect 1577 -337 1631 -336
rect 1835 -340 1839 -276
rect 1976 -323 1980 -259
rect 1998 -263 2003 -259
rect 2036 -262 2040 -259
rect 2087 -256 2092 -250
rect 2170 -256 2175 -250
rect 2087 -261 2175 -256
rect 2036 -267 2057 -262
rect 2013 -272 2018 -268
rect 1993 -277 2027 -272
rect 2021 -314 2026 -277
rect 2087 -284 2092 -261
rect 2136 -267 2139 -264
rect 2134 -272 2144 -267
rect 2042 -295 2047 -292
rect 2136 -284 2141 -272
rect 2053 -314 2058 -289
rect 2170 -284 2175 -261
rect 2184 -314 2189 -239
rect 2201 -277 2244 -272
rect 2203 -284 2208 -277
rect 2215 -284 2220 -277
rect 2230 -297 2235 -289
rect 2249 -297 2254 -217
rect 2215 -302 2218 -298
rect 2230 -302 2254 -297
rect 2230 -306 2235 -302
rect 2021 -315 2189 -314
rect 2215 -315 2220 -311
rect 2021 -319 2245 -315
rect 2184 -320 2245 -319
rect 1976 -328 2145 -323
rect 2140 -333 2145 -328
rect 2162 -333 2167 -329
rect 2140 -338 2167 -333
rect 1332 -350 1337 -345
rect 1310 -355 1337 -350
rect 1552 -349 1608 -344
rect 1366 -370 1372 -354
rect 1648 -350 1653 -346
rect 1670 -345 1839 -340
rect 1670 -350 1675 -345
rect 1648 -355 1675 -350
rect 1547 -368 1553 -365
rect 1706 -368 1711 -353
rect 1547 -371 1711 -368
rect 2108 -401 2245 -396
rect 2108 -403 2113 -401
rect 1980 -417 2085 -413
rect 1980 -418 2028 -417
rect 2004 -425 2009 -418
rect 2032 -429 2037 -417
rect 1989 -439 1994 -430
rect 2044 -429 2049 -417
rect 2127 -423 2180 -417
rect 2127 -429 2132 -423
rect 1967 -443 1994 -439
rect 2006 -443 2018 -439
rect 2023 -443 2031 -439
rect 1967 -507 1971 -443
rect 1989 -447 1994 -443
rect 2027 -446 2031 -443
rect 2078 -440 2083 -434
rect 2161 -440 2166 -434
rect 2078 -445 2166 -440
rect 2027 -451 2048 -446
rect 2004 -456 2009 -452
rect 1984 -461 2018 -456
rect 2012 -498 2017 -461
rect 2078 -468 2083 -445
rect 2127 -451 2130 -448
rect 2125 -456 2135 -451
rect 2033 -479 2038 -476
rect 2127 -468 2132 -456
rect 2044 -498 2049 -473
rect 2161 -468 2166 -445
rect 2175 -498 2180 -423
rect 2192 -461 2235 -456
rect 2194 -468 2199 -461
rect 2206 -468 2211 -461
rect 2221 -481 2226 -473
rect 2240 -481 2245 -401
rect 2206 -486 2209 -482
rect 2221 -486 2245 -481
rect 2221 -490 2226 -486
rect 2012 -499 2180 -498
rect 2206 -499 2211 -495
rect 2012 -503 2236 -499
rect 2175 -504 2236 -503
rect 1967 -512 2136 -507
rect 2131 -517 2136 -512
rect 2153 -517 2158 -513
rect 2131 -522 2158 -517
<< m2contact >>
rect 944 1020 949 1025
rect 895 1010 902 1017
rect 936 995 941 1002
rect 859 984 869 989
rect 944 984 950 989
rect 943 960 949 966
rect 882 929 889 936
rect 669 893 674 900
rect 866 897 872 906
rect 700 891 707 897
rect 795 880 800 886
rect 132 802 141 813
rect 655 864 661 869
rect 795 864 802 869
rect 1071 853 1086 862
rect 655 844 662 849
rect 795 844 802 849
rect 931 846 936 851
rect 186 777 199 787
rect 75 763 86 773
rect 461 761 475 771
rect 186 733 193 739
rect 229 708 234 713
rect 356 733 361 738
rect 227 690 232 695
rect 287 707 294 712
rect 250 690 255 695
rect 304 667 309 672
rect 383 695 390 702
rect 398 693 403 700
rect 458 690 463 695
rect 530 749 538 757
rect 604 823 615 830
rect 655 823 663 829
rect 736 824 750 829
rect 795 826 802 831
rect 578 701 587 715
rect 931 825 937 830
rect 840 789 853 805
rect 655 779 664 786
rect 681 777 690 785
rect 796 782 801 788
rect 899 789 909 798
rect 1077 792 1088 803
rect 1176 786 1187 795
rect 2362 822 2371 831
rect 2071 807 2083 818
rect 796 758 801 765
rect 615 743 622 748
rect 961 742 967 750
rect 1116 725 1126 731
rect 1206 717 1211 722
rect 1157 707 1164 714
rect 690 696 695 702
rect 706 696 711 702
rect 754 696 759 703
rect 472 665 477 670
rect 720 666 730 674
rect 755 672 765 680
rect 545 648 561 660
rect 503 599 517 608
rect 224 539 229 544
rect 183 510 190 516
rect 226 486 231 491
rect 353 511 358 516
rect 224 468 229 473
rect 286 482 292 488
rect 247 468 252 473
rect 379 473 388 478
rect 301 445 306 450
rect 455 468 460 473
rect 469 443 474 448
rect 568 647 585 658
rect 548 598 560 610
rect 621 623 633 634
rect 570 581 581 596
rect 541 558 552 569
rect 739 642 751 658
rect 914 629 925 638
rect 1198 692 1203 699
rect 1221 692 1226 699
rect 1012 623 1024 630
rect 1039 623 1051 630
rect 779 579 789 586
rect 815 577 828 587
rect 716 562 727 573
rect 958 560 970 574
rect 1102 568 1117 577
rect 1318 554 1326 561
rect 573 531 585 541
rect 651 532 662 541
rect 1663 762 1676 775
rect 1991 763 1998 771
rect 2618 794 2628 803
rect 2186 778 2194 785
rect 2114 770 2124 777
rect 2132 758 2142 766
rect 2262 774 2271 780
rect 2766 771 2776 781
rect 2281 759 2289 765
rect 1887 691 1892 696
rect 1980 698 1986 705
rect 1934 681 1941 688
rect 2023 691 2028 696
rect 2118 699 2124 706
rect 1872 666 1877 673
rect 1895 666 1900 673
rect 2070 681 2077 688
rect 2169 693 2174 698
rect 2264 700 2270 707
rect 2216 683 2223 690
rect 2316 693 2321 698
rect 2420 700 2427 708
rect 2008 666 2013 673
rect 2031 666 2036 673
rect 2154 668 2159 675
rect 2177 668 2182 675
rect 2363 683 2370 690
rect 2528 692 2533 697
rect 2281 667 2289 673
rect 2301 668 2306 675
rect 2324 668 2329 675
rect 2575 682 2582 689
rect 2664 692 2669 697
rect 2513 667 2518 674
rect 2536 667 2541 674
rect 2711 682 2718 689
rect 2810 694 2815 699
rect 2857 684 2864 691
rect 2957 694 2962 699
rect 2649 667 2654 674
rect 2672 667 2677 674
rect 2795 669 2800 676
rect 2818 669 2823 676
rect 3004 684 3011 691
rect 2942 669 2947 676
rect 2965 669 2970 676
rect 1887 583 1892 588
rect 1993 591 1998 597
rect 1934 573 1941 580
rect 2031 583 2036 588
rect 2133 589 2139 596
rect 1832 553 1838 560
rect 1872 557 1877 565
rect 1895 558 1900 565
rect 660 480 667 486
rect 759 471 764 476
rect 815 481 821 486
rect 710 461 717 468
rect 906 471 911 476
rect 959 478 966 484
rect 153 400 160 407
rect 198 401 205 408
rect 480 360 489 370
rect 144 348 152 354
rect 45 300 50 305
rect 161 326 168 332
rect 356 326 361 331
rect 228 299 233 305
rect 227 283 232 288
rect 147 267 153 273
rect 186 267 192 272
rect 226 255 231 261
rect 143 243 151 249
rect 288 298 293 303
rect 250 283 255 288
rect 304 260 309 265
rect 383 288 391 293
rect 458 283 463 288
rect 472 258 477 263
rect 542 432 554 443
rect 572 438 583 448
rect 751 446 756 453
rect 774 446 779 453
rect 857 461 864 468
rect 1052 469 1057 474
rect 1103 476 1109 481
rect 898 446 903 453
rect 1003 459 1010 466
rect 1188 469 1193 474
rect 921 446 926 453
rect 1044 444 1049 451
rect 1067 444 1072 451
rect 1139 459 1146 466
rect 1180 444 1185 451
rect 1203 444 1208 451
rect 541 376 551 389
rect 535 349 545 357
rect 635 373 641 378
rect 620 324 630 334
rect 501 225 510 232
rect 502 196 509 203
rect 510 168 516 176
rect 186 151 193 157
rect 356 151 361 156
rect 228 125 233 130
rect 227 108 232 113
rect 288 123 294 128
rect 250 108 255 113
rect 378 113 388 118
rect 304 85 309 90
rect 458 108 463 113
rect 472 83 477 88
rect 617 95 626 107
rect 476 38 485 48
rect 1580 513 1585 518
rect 1660 522 1666 527
rect 2078 573 2085 580
rect 2180 585 2185 590
rect 2282 592 2288 598
rect 2227 575 2234 582
rect 2325 586 2330 591
rect 2407 592 2415 599
rect 2372 576 2379 583
rect 2016 558 2021 565
rect 2039 558 2044 565
rect 2165 560 2170 567
rect 2188 560 2193 567
rect 2310 560 2315 567
rect 2333 561 2338 568
rect 1627 504 1634 510
rect 1488 482 1496 490
rect 1565 489 1570 496
rect 1656 501 1665 510
rect 1832 518 1838 523
rect 1588 490 1593 496
rect 662 371 668 377
rect 750 364 755 369
rect 804 373 809 378
rect 701 354 708 361
rect 895 363 900 368
rect 945 369 952 374
rect 742 339 747 346
rect 765 338 770 345
rect 846 353 853 360
rect 1044 361 1049 366
rect 1090 370 1095 375
rect 1405 383 1410 388
rect 1429 383 1435 388
rect 1442 383 1447 388
rect 1465 383 1473 388
rect 887 338 892 345
rect 910 338 915 345
rect 995 351 1002 358
rect 1188 361 1193 366
rect 1337 363 1353 375
rect 1036 336 1041 343
rect 1059 336 1064 343
rect 1139 351 1146 358
rect 1180 336 1185 343
rect 1203 335 1208 343
rect 1244 335 1249 341
rect 1318 335 1323 341
rect 1441 361 1447 366
rect 1319 171 1326 177
rect 1720 503 1729 512
rect 1791 485 1796 490
rect 1666 404 1671 409
rect 1579 395 1584 400
rect 1624 386 1632 391
rect 1564 370 1569 375
rect 1586 369 1592 375
rect 1848 475 1855 484
rect 2383 460 2388 465
rect 1732 404 1738 409
rect 2218 394 2223 399
rect 2288 403 2293 408
rect 2335 393 2342 400
rect 2424 403 2429 408
rect 2273 378 2278 385
rect 2296 378 2301 385
rect 1762 361 1769 369
rect 2099 351 2104 356
rect 2471 393 2478 400
rect 2570 405 2575 410
rect 2617 395 2624 402
rect 2717 405 2722 410
rect 2409 378 2414 385
rect 2432 378 2437 385
rect 2555 380 2560 387
rect 2578 380 2583 387
rect 2764 395 2771 402
rect 2702 380 2707 387
rect 2725 380 2730 387
rect 1670 300 1678 306
rect 1578 291 1583 296
rect 1623 282 1631 288
rect 2002 228 2007 233
rect 1578 195 1583 200
rect 1805 203 1815 210
rect 1624 185 1632 191
rect 1769 185 1774 190
rect 1586 171 1591 178
rect 1938 184 1944 189
rect 2006 156 2011 161
rect 2288 295 2293 300
rect 2367 304 2372 309
rect 2335 285 2342 292
rect 2520 304 2525 309
rect 2432 295 2437 300
rect 2273 269 2278 277
rect 2296 270 2301 277
rect 2479 285 2486 292
rect 2667 306 2674 311
rect 2581 297 2586 302
rect 2628 287 2635 294
rect 2812 307 2819 312
rect 2726 298 2731 303
rect 2773 288 2780 295
rect 2417 270 2422 277
rect 2440 270 2445 277
rect 2566 272 2571 279
rect 2589 272 2594 279
rect 2711 272 2716 279
rect 2734 273 2739 280
rect 1831 123 1839 136
rect 2036 122 2042 127
rect 671 92 685 107
rect 2112 121 2117 126
rect 288 0 299 11
rect 2046 95 2051 100
rect 2006 78 2012 84
rect 2147 83 2152 88
rect 2060 55 2065 60
rect 2214 78 2219 83
rect 2228 53 2233 58
rect 1579 -47 1585 -40
rect 1539 -61 1544 -56
rect 1555 -62 1560 -57
rect 1571 -62 1576 -57
rect 2106 -62 2111 -57
rect 2038 -87 2043 -82
rect 1230 -208 1239 -202
rect 1271 -144 1276 -139
rect 1368 -152 1373 -147
rect 1418 -145 1423 -140
rect 1319 -162 1326 -155
rect 1514 -154 1519 -149
rect 1559 -145 1564 -140
rect 1360 -177 1365 -170
rect 1465 -164 1472 -157
rect 1650 -154 1655 -149
rect 1383 -177 1388 -170
rect 1278 -188 1290 -181
rect 1506 -179 1511 -172
rect 1529 -179 1534 -172
rect 1601 -164 1608 -157
rect 1642 -179 1647 -172
rect 1665 -179 1670 -172
rect 1439 -198 1446 -193
rect 1280 -208 1289 -201
rect 1642 -198 1647 -191
rect 1785 -196 1792 -189
rect 1727 -205 1734 -200
rect 1258 -225 1271 -217
rect 1439 -238 1446 -230
rect 1378 -251 1383 -246
rect 1276 -294 1281 -289
rect 1262 -319 1267 -314
rect 1229 -340 1236 -331
rect 1366 -278 1372 -272
rect 1343 -289 1348 -284
rect 1441 -277 1446 -272
rect 1430 -317 1435 -312
rect 1451 -337 1458 -331
rect 1999 -105 2004 -100
rect 2141 -100 2146 -95
rect 2054 -128 2059 -123
rect 2208 -105 2213 -100
rect 2222 -130 2227 -125
rect 1716 -251 1721 -246
rect 1614 -294 1619 -289
rect 1600 -319 1605 -314
rect 1570 -337 1577 -331
rect 2094 -234 2099 -229
rect 2027 -259 2032 -254
rect 1706 -278 1711 -273
rect 1681 -289 1686 -284
rect 1779 -277 1784 -272
rect 1768 -317 1773 -312
rect 1988 -278 1993 -272
rect 2129 -272 2134 -267
rect 2042 -300 2047 -295
rect 2196 -277 2201 -272
rect 2210 -302 2215 -297
rect 1366 -354 1372 -348
rect 1608 -349 1615 -343
rect 1706 -353 1711 -348
rect 1547 -365 1554 -357
rect 2085 -418 2090 -413
rect 2018 -443 2023 -438
rect 1979 -462 1984 -455
rect 2120 -456 2125 -451
rect 2033 -484 2038 -479
rect 2187 -461 2192 -456
rect 2201 -486 2206 -481
<< metal2 >>
rect 918 1020 944 1023
rect 918 1016 923 1020
rect 902 1011 923 1016
rect 632 995 936 998
rect 632 993 941 995
rect 633 914 636 993
rect 869 984 888 989
rect 883 936 888 984
rect 944 966 947 984
rect 46 911 636 914
rect 46 761 50 911
rect 655 893 669 895
rect 872 899 906 904
rect 655 891 674 893
rect 707 892 824 895
rect 754 891 824 892
rect 655 869 659 891
rect 796 869 800 880
rect 342 856 1071 860
rect 125 804 132 809
rect 343 788 348 856
rect 554 825 604 829
rect 655 829 660 844
rect 742 829 746 856
rect 796 831 800 844
rect 931 830 935 846
rect 1925 843 1932 844
rect 1925 842 2193 843
rect 1925 838 2194 842
rect 571 815 1257 819
rect 199 777 283 785
rect 178 769 234 770
rect 86 767 234 769
rect 343 767 349 788
rect 86 764 349 767
rect 86 763 184 764
rect 45 680 50 761
rect 45 305 49 680
rect 154 407 158 740
rect 186 516 189 733
rect 229 713 234 764
rect 364 761 461 767
rect 364 758 471 761
rect 364 738 369 758
rect 361 733 383 738
rect 232 690 250 695
rect 288 590 293 707
rect 377 695 383 733
rect 390 695 398 700
rect 458 695 463 758
rect 571 754 580 815
rect 731 798 840 799
rect 645 793 840 798
rect 645 792 759 793
rect 538 749 580 754
rect 615 779 655 784
rect 681 785 688 792
rect 853 793 856 799
rect 1008 794 1077 797
rect 909 792 1077 794
rect 909 789 1081 792
rect 615 748 621 779
rect 796 765 800 782
rect 961 750 966 778
rect 1116 731 1120 792
rect 1177 720 1182 786
rect 1251 774 1257 815
rect 1925 809 1932 838
rect 1612 803 1932 809
rect 1955 817 1960 818
rect 1955 811 2071 817
rect 1177 717 1206 720
rect 556 706 578 712
rect 304 625 309 667
rect 462 665 472 669
rect 462 625 468 665
rect 556 660 562 706
rect 1177 713 1185 717
rect 1164 708 1185 713
rect 1250 697 1257 774
rect 1226 694 1257 697
rect 1226 693 1254 694
rect 1198 688 1203 692
rect 714 666 720 672
rect 561 648 562 660
rect 585 647 739 655
rect 304 624 610 625
rect 304 620 612 624
rect 633 629 720 630
rect 633 623 721 629
rect 457 619 612 620
rect 596 617 612 619
rect 517 599 548 606
rect 288 585 570 590
rect 186 359 189 510
rect 226 491 229 539
rect 361 536 468 545
rect 361 516 366 536
rect 358 511 380 516
rect 229 468 247 473
rect 205 402 232 406
rect 161 355 189 359
rect 161 354 164 355
rect 152 348 164 354
rect 228 352 232 402
rect 287 383 291 482
rect 374 478 380 511
rect 374 473 379 478
rect 455 473 460 536
rect 301 403 306 445
rect 459 443 469 447
rect 542 443 548 558
rect 575 448 580 531
rect 459 403 465 443
rect 301 400 465 403
rect 301 398 565 400
rect 454 397 565 398
rect 287 379 541 383
rect 398 364 480 368
rect 161 332 164 348
rect 200 349 232 352
rect 200 337 205 349
rect 186 334 205 337
rect 146 267 147 272
rect 146 249 149 267
rect 161 249 164 326
rect 186 272 190 334
rect 228 305 232 349
rect 364 351 471 360
rect 364 331 369 351
rect 361 326 383 331
rect 232 283 250 288
rect 161 245 189 249
rect 186 157 189 245
rect 228 130 231 255
rect 289 200 293 298
rect 377 288 383 326
rect 458 288 463 351
rect 304 218 309 260
rect 462 258 472 262
rect 462 218 468 258
rect 537 230 542 349
rect 560 328 565 397
rect 510 227 542 230
rect 510 226 541 227
rect 304 216 468 218
rect 558 217 565 328
rect 600 290 610 617
rect 634 591 640 592
rect 634 586 706 591
rect 634 488 640 586
rect 699 557 705 586
rect 716 573 721 623
rect 758 557 763 672
rect 1613 662 1621 803
rect 1955 789 1960 811
rect 2188 816 2194 838
rect 2362 831 3074 835
rect 2371 827 3074 831
rect 802 652 1621 662
rect 781 563 787 579
rect 699 553 763 557
rect 780 539 787 563
rect 662 532 787 539
rect 620 487 656 488
rect 620 486 664 487
rect 620 482 660 486
rect 620 334 628 482
rect 633 481 660 482
rect 733 471 759 474
rect 733 467 738 471
rect 717 462 738 467
rect 803 451 810 652
rect 1613 651 1621 652
rect 1635 781 1960 789
rect 1979 785 2156 790
rect 2188 785 2193 816
rect 2628 794 2629 803
rect 2246 785 2456 790
rect 1979 784 2006 785
rect 1635 641 1641 781
rect 943 634 1642 641
rect 815 555 819 577
rect 918 555 923 629
rect 815 551 924 555
rect 815 486 819 551
rect 880 471 906 474
rect 880 467 885 471
rect 864 462 885 467
rect 779 448 810 451
rect 779 447 807 448
rect 751 428 756 446
rect 898 428 903 446
rect 943 450 950 634
rect 1007 623 1012 629
rect 1024 623 1039 630
rect 959 554 963 560
rect 1007 554 1014 623
rect 1664 612 1670 762
rect 1980 705 1986 784
rect 2118 777 2123 778
rect 1892 691 1918 694
rect 1913 687 1918 691
rect 1913 682 1934 687
rect 1092 607 1670 612
rect 1772 661 1777 663
rect 1872 662 1877 666
rect 1855 661 1877 662
rect 1772 657 1877 661
rect 1772 656 1861 657
rect 1092 604 1731 607
rect 959 548 1015 554
rect 959 484 963 548
rect 1026 469 1052 472
rect 1026 465 1031 469
rect 1010 460 1031 465
rect 926 446 950 450
rect 921 445 948 446
rect 1092 447 1097 604
rect 1733 603 1737 604
rect 1253 590 1260 591
rect 1772 590 1777 656
rect 1253 584 1777 590
rect 1103 563 1109 568
rect 1103 557 1199 563
rect 1103 481 1109 557
rect 1162 469 1188 472
rect 1162 465 1167 469
rect 1146 460 1167 465
rect 1072 444 1098 447
rect 1044 428 1049 444
rect 1180 428 1185 444
rect 1253 446 1260 584
rect 1772 582 1777 584
rect 1208 444 1260 446
rect 1203 441 1260 444
rect 1318 500 1323 554
rect 1666 523 1768 527
rect 1585 513 1611 516
rect 1606 509 1611 513
rect 1606 505 1627 509
rect 1606 504 1618 505
rect 751 425 1270 428
rect 641 373 662 377
rect 724 364 750 367
rect 804 368 807 373
rect 724 360 729 364
rect 869 363 895 366
rect 708 355 729 360
rect 869 359 874 363
rect 853 354 874 359
rect 945 361 948 369
rect 1018 361 1044 364
rect 1018 357 1023 361
rect 1002 352 1023 357
rect 1090 350 1094 370
rect 1162 361 1188 364
rect 1162 357 1167 361
rect 1146 352 1167 357
rect 742 314 747 339
rect 770 339 792 343
rect 887 314 892 338
rect 915 338 931 340
rect 910 336 931 338
rect 1064 336 1074 340
rect 1036 314 1041 336
rect 1180 314 1185 336
rect 1208 335 1244 339
rect 1266 314 1270 425
rect 1318 371 1324 500
rect 1433 482 1488 487
rect 1565 487 1570 489
rect 1496 482 1570 487
rect 1433 390 1438 482
rect 1588 472 1593 490
rect 1520 465 1593 472
rect 1433 388 1437 390
rect 1520 388 1527 465
rect 1584 395 1607 398
rect 1388 383 1405 388
rect 1435 383 1437 388
rect 1473 383 1527 388
rect 1602 391 1607 395
rect 1611 391 1616 504
rect 1665 504 1720 510
rect 1671 404 1732 409
rect 1602 386 1624 391
rect 1318 364 1337 371
rect 1388 357 1394 383
rect 1442 366 1446 383
rect 1520 371 1527 383
rect 1520 370 1564 371
rect 1520 364 1569 370
rect 1586 357 1592 369
rect 1388 353 1592 357
rect 1388 352 1394 353
rect 742 311 1270 314
rect 742 310 747 311
rect 600 287 1090 290
rect 600 286 610 287
rect 896 266 900 271
rect 895 263 946 266
rect 953 263 954 266
rect 895 262 954 263
rect 772 248 805 251
rect 772 247 810 248
rect 558 216 616 217
rect 896 216 900 262
rect 1080 232 1247 238
rect 304 213 551 216
rect 289 196 502 200
rect 364 176 471 185
rect 510 176 516 182
rect 364 156 369 176
rect 361 151 383 156
rect 232 108 250 113
rect 288 28 292 123
rect 377 118 383 151
rect 377 113 378 118
rect 458 113 463 176
rect 304 43 309 85
rect 462 83 472 87
rect 462 44 468 83
rect 461 43 476 44
rect 304 38 476 43
rect 542 42 551 213
rect 558 213 903 216
rect 558 210 616 213
rect 940 216 1218 218
rect 940 212 1219 216
rect 800 184 1182 188
rect 626 95 671 104
rect 749 44 759 45
rect 631 43 759 44
rect 571 42 759 43
rect 542 39 759 42
rect 542 38 749 39
rect 1177 48 1182 184
rect 1209 81 1219 212
rect 1242 211 1247 232
rect 1242 133 1248 211
rect 1266 150 1270 311
rect 1319 177 1322 335
rect 1428 171 1432 353
rect 1583 291 1607 294
rect 1602 287 1607 291
rect 1611 287 1616 386
rect 1719 351 1722 404
rect 1763 369 1768 523
rect 1792 490 1795 656
rect 1895 650 1900 666
rect 1991 670 1996 763
rect 2118 706 2123 770
rect 2151 758 2156 785
rect 2246 758 2250 785
rect 2028 691 2054 694
rect 2049 687 2054 691
rect 2049 682 2070 687
rect 1991 666 2008 670
rect 2134 671 2139 758
rect 2151 754 2250 758
rect 2264 707 2269 774
rect 2281 755 2285 759
rect 2281 752 2402 755
rect 2174 693 2200 696
rect 2195 689 2200 693
rect 2195 684 2216 689
rect 2134 668 2154 671
rect 2134 667 2159 668
rect 2139 666 2155 667
rect 1991 665 2005 666
rect 1991 664 1996 665
rect 2031 650 2036 666
rect 2177 650 2182 668
rect 2281 673 2285 752
rect 2421 708 2427 755
rect 2321 693 2347 696
rect 2342 689 2347 693
rect 2342 684 2363 689
rect 2289 671 2297 672
rect 2289 668 2301 671
rect 2289 667 2306 668
rect 2324 650 2329 668
rect 2450 662 2456 785
rect 2533 692 2559 695
rect 2554 688 2559 692
rect 2554 683 2575 688
rect 2513 662 2518 667
rect 2450 657 2518 662
rect 2625 671 2629 794
rect 2776 771 2777 780
rect 2669 692 2695 695
rect 2690 688 2695 692
rect 2690 683 2711 688
rect 2624 667 2649 671
rect 2771 673 2777 771
rect 2915 753 2916 760
rect 2815 694 2841 697
rect 2836 690 2841 694
rect 2836 685 2857 690
rect 2771 672 2789 673
rect 2771 669 2795 672
rect 2771 668 2800 669
rect 2911 672 2916 753
rect 2962 694 2988 697
rect 2983 690 2988 694
rect 2983 685 3004 690
rect 1810 647 2329 650
rect 1810 536 1814 647
rect 1892 583 1918 586
rect 1913 579 1918 583
rect 1993 580 1998 591
rect 2415 594 2456 599
rect 2036 583 2062 586
rect 1913 574 1934 579
rect 2057 579 2062 583
rect 2057 574 2078 579
rect 2133 568 2139 589
rect 2185 585 2211 588
rect 2206 581 2211 585
rect 2206 576 2227 581
rect 2284 570 2288 592
rect 2330 586 2356 589
rect 2351 582 2356 586
rect 2351 577 2372 582
rect 1861 560 1872 561
rect 1838 557 1872 560
rect 1895 536 1900 558
rect 2010 558 2016 561
rect 2010 557 2021 558
rect 2039 536 2044 558
rect 2159 560 2165 563
rect 2159 559 2170 560
rect 2188 536 2193 560
rect 2306 560 2310 564
rect 2333 536 2338 561
rect 1810 533 2338 536
rect 1810 526 1814 533
rect 2333 532 2338 533
rect 1806 523 1814 526
rect 1719 348 1772 351
rect 1669 300 1670 304
rect 1678 300 1719 304
rect 1602 282 1623 287
rect 1583 195 1606 198
rect 1602 191 1606 195
rect 1611 191 1616 282
rect 1602 186 1624 191
rect 1428 168 1591 171
rect 1586 167 1591 168
rect 1713 150 1719 300
rect 1769 190 1772 348
rect 1806 210 1810 523
rect 2154 522 2158 523
rect 1834 495 1837 518
rect 1833 314 1837 495
rect 1848 484 1854 490
rect 2006 458 2010 493
rect 2154 468 2158 516
rect 2364 471 2367 526
rect 2536 490 2541 667
rect 2672 505 2677 667
rect 2818 521 2823 669
rect 2910 669 2942 672
rect 2910 668 2947 669
rect 2965 651 2970 669
rect 2966 602 2970 651
rect 3067 474 3074 827
rect 1892 449 2010 458
rect 2153 459 2158 468
rect 2177 466 2367 471
rect 2528 467 3074 474
rect 1266 145 1719 150
rect 1713 144 1719 145
rect 1833 136 1837 308
rect 1892 284 1897 449
rect 1919 419 1928 421
rect 2153 419 2157 459
rect 1919 411 2160 419
rect 1243 105 1248 133
rect 1892 105 1897 276
rect 1919 228 1928 411
rect 2177 397 2189 466
rect 2293 403 2319 406
rect 2314 399 2319 403
rect 1966 385 2189 397
rect 2223 394 2258 397
rect 2314 394 2335 399
rect 1926 218 1928 228
rect 1243 99 1902 105
rect 1209 76 1218 81
rect 1919 76 1928 218
rect 1967 191 1977 385
rect 2255 381 2258 394
rect 2255 378 2273 381
rect 2383 381 2386 460
rect 2429 403 2455 406
rect 2450 399 2455 403
rect 2450 394 2471 399
rect 2383 378 2409 381
rect 2529 384 2534 467
rect 2575 405 2601 408
rect 2596 401 2601 405
rect 2596 396 2617 401
rect 2529 380 2555 384
rect 2681 383 2685 407
rect 2722 405 2748 408
rect 2743 401 2748 405
rect 2743 396 2764 401
rect 2681 380 2702 383
rect 2296 362 2301 378
rect 2432 362 2437 378
rect 2578 362 2583 380
rect 2725 362 2730 380
rect 2211 359 2730 362
rect 2211 354 2215 359
rect 2104 351 2215 354
rect 2211 248 2215 351
rect 2372 304 2379 309
rect 2525 304 2534 308
rect 2674 306 2683 310
rect 2819 303 2822 312
rect 2293 295 2319 298
rect 2437 295 2463 298
rect 2586 297 2612 300
rect 2731 298 2757 301
rect 2314 291 2319 295
rect 2251 275 2254 291
rect 2314 286 2335 291
rect 2458 291 2463 295
rect 2607 293 2612 297
rect 2752 294 2757 298
rect 2458 286 2479 291
rect 2607 288 2628 293
rect 2752 289 2773 294
rect 2251 271 2273 275
rect 2296 248 2301 270
rect 2404 270 2417 274
rect 2422 270 2423 274
rect 2404 269 2423 270
rect 2552 272 2566 276
rect 2552 271 2571 272
rect 2690 273 2711 277
rect 2440 248 2445 270
rect 2589 248 2594 272
rect 2734 248 2739 273
rect 2211 245 2739 248
rect 2734 244 2739 245
rect 2007 228 2042 233
rect 1939 177 1943 184
rect 1209 66 1930 76
rect 1938 70 1943 177
rect 1919 64 1928 66
rect 1967 48 1977 183
rect 1177 39 1977 48
rect 2006 84 2010 156
rect 2036 127 2041 228
rect 2120 154 2227 155
rect 2120 151 2297 154
rect 2120 146 2227 151
rect 2120 126 2125 146
rect 2117 121 2139 126
rect 288 11 293 28
rect 2006 -7 2011 78
rect 1999 -12 2011 -7
rect 2046 70 2051 95
rect 2133 88 2139 121
rect 2133 83 2147 88
rect 2214 83 2219 146
rect 2046 64 2047 70
rect 2139 69 2144 83
rect 1579 -40 1625 -39
rect 1585 -44 1625 -40
rect 1273 -60 1539 -57
rect 1273 -139 1276 -60
rect 1555 -66 1560 -62
rect 1538 -70 1560 -66
rect 1538 -81 1542 -70
rect 1571 -74 1576 -62
rect 1419 -86 1542 -81
rect 1559 -79 1576 -74
rect 1419 -140 1423 -86
rect 1559 -140 1563 -79
rect 1342 -152 1368 -149
rect 1342 -156 1347 -152
rect 1326 -161 1347 -156
rect 1488 -154 1514 -151
rect 1619 -151 1625 -44
rect 1619 -154 1650 -151
rect 1488 -158 1493 -154
rect 1472 -163 1493 -158
rect 1619 -158 1629 -154
rect 1608 -163 1629 -158
rect 1210 -188 1278 -183
rect 1211 -331 1215 -188
rect 1239 -208 1280 -202
rect 1360 -202 1365 -177
rect 1383 -194 1388 -177
rect 1383 -198 1439 -194
rect 1506 -194 1511 -179
rect 1446 -198 1511 -194
rect 1529 -194 1534 -179
rect 1642 -191 1647 -179
rect 1529 -198 1642 -194
rect 1665 -200 1670 -179
rect 1727 -200 1734 -55
rect 1786 -189 1792 -56
rect 1999 -100 2004 -12
rect 2046 -52 2051 64
rect 2060 13 2065 55
rect 2218 53 2228 57
rect 2218 52 2232 53
rect 2218 16 2224 52
rect 2060 8 2216 13
rect 1665 -202 1727 -200
rect 1360 -205 1727 -202
rect 1734 -205 1784 -200
rect 1271 -225 1713 -217
rect 1268 -226 1713 -225
rect 1276 -289 1281 -226
rect 1370 -246 1375 -226
rect 1356 -251 1378 -246
rect 1356 -284 1362 -251
rect 1441 -272 1446 -238
rect 1348 -289 1362 -284
rect 1351 -303 1356 -289
rect 1267 -319 1277 -315
rect 1211 -337 1229 -331
rect 1271 -359 1277 -319
rect 1366 -348 1372 -278
rect 1614 -289 1619 -226
rect 1708 -246 1713 -226
rect 1694 -251 1716 -246
rect 1694 -284 1700 -251
rect 1779 -272 1784 -205
rect 1999 -221 2004 -105
rect 2038 -55 2051 -52
rect 2114 -33 2221 -28
rect 2293 -33 2296 151
rect 2114 -36 2297 -33
rect 2114 -37 2221 -36
rect 2038 -82 2043 -55
rect 2114 -57 2119 -37
rect 2111 -62 2133 -57
rect 2038 -169 2043 -87
rect 2127 -95 2133 -62
rect 2127 -100 2141 -95
rect 2208 -100 2213 -37
rect 2133 -114 2138 -100
rect 1686 -289 1700 -284
rect 1988 -225 2004 -221
rect 2027 -173 2043 -169
rect 2054 -170 2059 -128
rect 2212 -130 2222 -126
rect 2212 -131 2226 -130
rect 2212 -167 2218 -131
rect 1988 -272 1992 -225
rect 2027 -254 2032 -173
rect 2054 -175 2211 -170
rect 2102 -201 2209 -200
rect 2293 -201 2296 -36
rect 2102 -205 2296 -201
rect 2102 -209 2209 -205
rect 2102 -229 2107 -209
rect 2099 -234 2121 -229
rect 1689 -303 1694 -289
rect 1430 -358 1435 -317
rect 1605 -319 1615 -315
rect 1458 -337 1570 -331
rect 1609 -343 1615 -319
rect 1430 -359 1547 -358
rect 1271 -363 1547 -359
rect 1271 -364 1435 -363
rect 1609 -359 1615 -349
rect 1706 -348 1711 -278
rect 1768 -359 1773 -317
rect 1609 -364 1773 -359
rect 1988 -399 1992 -278
rect 2027 -345 2032 -259
rect 2115 -267 2121 -234
rect 2115 -272 2129 -267
rect 2196 -272 2201 -209
rect 2121 -286 2126 -272
rect 1979 -403 1992 -399
rect 2018 -348 2032 -345
rect 2042 -342 2047 -300
rect 2200 -302 2210 -298
rect 2200 -303 2214 -302
rect 2200 -340 2206 -303
rect 2042 -347 2199 -342
rect 1979 -455 1983 -403
rect 2018 -438 2022 -348
rect 2293 -374 2296 -205
rect 2291 -383 2296 -374
rect 2189 -384 2296 -383
rect 2093 -388 2296 -384
rect 2093 -393 2200 -388
rect 2093 -413 2098 -393
rect 2090 -418 2112 -413
rect 2106 -451 2112 -418
rect 2106 -456 2120 -451
rect 2187 -456 2192 -393
rect 2112 -470 2117 -456
rect 2033 -526 2038 -484
rect 2191 -486 2201 -482
rect 2191 -487 2205 -486
rect 2191 -524 2197 -487
rect 2033 -531 2191 -526
rect 2186 -532 2191 -531
<< m3contact >>
rect 906 898 913 904
rect 824 888 837 896
rect 113 801 125 813
rect 546 824 554 833
rect 283 776 299 788
rect 152 740 160 748
rect 631 790 645 801
rect 1114 792 1127 799
rect 959 778 967 783
rect 1197 682 1205 688
rect 706 666 714 674
rect 387 364 398 372
rect 1731 604 1737 609
rect 1199 557 1207 563
rect 804 363 809 368
rect 945 356 950 361
rect 1090 345 1095 350
rect 792 339 797 345
rect 931 335 938 341
rect 1074 336 1080 343
rect 1090 286 1095 291
rect 946 263 953 269
rect 763 246 772 254
rect 805 248 812 254
rect 1072 232 1080 242
rect 510 182 517 190
rect 931 212 940 221
rect 795 184 800 192
rect 759 36 771 49
rect 2402 752 2407 758
rect 2421 755 2429 763
rect 2906 753 2915 763
rect 2456 592 2466 600
rect 1993 574 1998 580
rect 2004 555 2010 563
rect 2132 561 2139 568
rect 2153 556 2159 564
rect 2283 563 2289 570
rect 2298 558 2306 568
rect 2361 526 2368 532
rect 2153 516 2160 522
rect 1848 490 1855 497
rect 2004 493 2012 500
rect 2965 593 2975 602
rect 2816 513 2826 521
rect 2669 498 2679 505
rect 2536 482 2543 490
rect 1833 308 1839 314
rect 1891 276 1898 284
rect 1917 218 1926 228
rect 2681 407 2686 412
rect 2379 304 2385 309
rect 2534 304 2539 309
rect 2683 306 2688 311
rect 2251 291 2256 296
rect 2817 298 2822 303
rect 2397 269 2404 274
rect 2547 271 2552 276
rect 2684 273 2690 278
rect 1966 183 1977 191
rect 1938 64 1945 70
rect 2047 64 2053 70
rect 2216 8 2224 16
rect 2211 -175 2218 -167
rect 2199 -348 2207 -340
rect 2191 -532 2199 -524
<< metal3 >>
rect 913 898 1033 903
rect 1029 889 1033 898
rect 829 886 1000 888
rect 1029 886 1119 889
rect 829 884 1001 886
rect 1029 884 1121 886
rect 154 831 157 832
rect 152 826 546 831
rect 116 393 120 801
rect 154 748 157 826
rect 390 797 394 799
rect 535 797 631 798
rect 389 793 631 797
rect 390 785 394 793
rect 535 791 631 793
rect 299 776 395 785
rect 997 783 1001 884
rect 1116 799 1121 884
rect 2402 841 3087 845
rect 967 778 1002 783
rect 2402 758 2406 841
rect 2429 761 2439 762
rect 2429 756 2906 761
rect 2429 755 2439 756
rect 607 601 615 603
rect 707 601 712 666
rect 606 594 713 601
rect 580 410 587 412
rect 607 410 615 594
rect 1199 563 1202 682
rect 1733 563 1737 604
rect 2461 600 2965 602
rect 2466 593 2965 600
rect 1781 567 1852 570
rect 1781 563 1785 567
rect 1733 559 1785 563
rect 1848 497 1852 567
rect 1993 485 1998 574
rect 2005 500 2010 555
rect 2132 505 2139 561
rect 2154 522 2158 556
rect 2283 518 2289 563
rect 2300 530 2303 558
rect 2300 527 2361 530
rect 2283 513 2816 518
rect 2132 499 2669 505
rect 1993 482 2536 485
rect 3081 486 3087 841
rect 2673 482 3087 486
rect 1993 481 2542 482
rect 2673 412 2676 482
rect 580 403 616 410
rect 2673 408 2681 412
rect 116 389 248 393
rect 240 369 245 389
rect 240 365 387 369
rect 580 292 587 403
rect 797 339 798 344
rect 579 188 587 292
rect 517 182 587 188
rect 761 246 763 252
rect 761 49 766 246
rect 795 192 798 339
rect 806 254 809 363
rect 931 221 937 335
rect 946 269 949 356
rect 1073 336 1074 338
rect 1073 242 1079 336
rect 1090 291 1094 345
rect 1839 308 2254 312
rect 2251 296 2254 308
rect 2381 296 2385 304
rect 2534 294 2538 304
rect 2684 298 2688 306
rect 2819 289 2822 298
rect 1898 276 2188 281
rect 2182 237 2188 276
rect 2399 237 2404 269
rect 2182 231 2404 237
rect 2547 224 2552 271
rect 1926 218 2552 224
rect 2684 191 2689 273
rect 1977 183 2689 191
rect 1945 64 2047 70
rect 2224 8 2379 13
rect 2218 -175 2402 -170
rect 2207 -346 2418 -341
rect 2199 -531 2444 -527
<< m4contact >>
rect 2381 291 2386 296
rect 2534 289 2539 294
rect 2683 293 2689 298
rect 2818 284 2823 289
rect 2379 8 2384 13
rect 2402 -175 2408 -168
rect 2418 -347 2426 -340
rect 2444 -533 2450 -525
<< metal4 >>
rect 2381 13 2384 291
rect 2685 289 2689 293
rect 2402 162 2407 163
rect 2534 162 2538 289
rect 2685 286 2699 289
rect 2694 171 2699 286
rect 2820 245 2823 284
rect 2750 244 2823 245
rect 2749 241 2823 244
rect 2749 233 2753 241
rect 2820 240 2823 241
rect 2402 158 2538 162
rect 2549 166 2699 171
rect 2707 229 2754 233
rect 2402 -168 2407 158
rect 2549 144 2554 166
rect 2707 152 2710 229
rect 2419 140 2554 144
rect 2572 148 2710 152
rect 2419 139 2553 140
rect 2419 -340 2424 139
rect 2572 126 2575 148
rect 2445 122 2575 126
rect 2445 -525 2449 122
<< labels >>
rlabel metal1 1426 386 1426 386 1 S0c
rlabel metal1 1411 386 1411 386 1 S0
rlabel metal1 1449 387 1449 387 1 S1
rlabel metal1 1665 406 1665 406 1 D1
rlabel metal1 1659 525 1659 525 1 D0
rlabel metal1 1667 206 1667 206 1 D3
rlabel metal1 1576 189 1576 189 1 DEC_AND_NODE_4
rlabel metal1 1576 212 1576 212 1 DEC_D3_NAND
rlabel metal1 1668 302 1668 302 1 D2
rlabel metal1 1577 285 1577 285 1 DEC_AND_NODE_3
rlabel metal1 1577 308 1577 308 1 DEC_D2_NAND
rlabel metal1 1579 389 1579 389 1 Dec_AND_node_2
rlabel metal1 1580 412 1580 412 1 DEC_D1_NAND
rlabel metal1 1575 531 1575 531 1 DEC_D0_NAND
rlabel metal1 1580 508 1580 508 1 Dec_AND_node_1
rlabel m2contact 1468 386 1468 386 1 S1c
rlabel metal1 1468 368 1468 368 1 gnd
rlabel metal1 1444 412 1444 412 1 vdd
rlabel metal2 1867 559 1867 559 1 B3
rlabel m3contact 2008 560 2008 560 1 B2
rlabel metal2 2160 562 2160 562 1 B1
rlabel metal1 2326 580 2326 580 1 ander_node_5
rlabel metal1 2178 580 2178 580 1 ander_node_6
rlabel metal1 2029 576 2029 576 1 ander_node_7
rlabel metal1 1884 578 1884 578 1 ander_node_8
rlabel metal1 2360 597 2360 597 1 and_b0e_nand
rlabel metal1 2225 596 2225 596 1 and_b1e_nand
rlabel metal1 2071 593 2071 593 1 and_b2e_nand
rlabel metal1 1923 593 1923 593 1 and_b3e_nand
rlabel metal1 2404 597 2404 597 1 and_b0e
rlabel metal1 2260 596 2260 596 1 and_b1e
rlabel metal1 2112 593 2112 593 1 and_b2e
rlabel metal1 1968 594 1968 594 1 and_b3e
rlabel metal1 2395 703 2395 703 1 and_a0e
rlabel metal1 2248 703 2248 703 1 and_a1e
rlabel metal1 2101 701 2101 701 1 and_a2e
rlabel metal1 1966 702 1966 702 1 and_a3e
rlabel metal1 2358 703 2358 703 1 and_a0e_nand
rlabel metal1 2212 704 2212 704 1 and_a1e_nand
rlabel metal1 2069 702 2069 702 1 and_a2e_nand
rlabel metal1 1925 703 1925 703 1 and_a3e_nand
rlabel metal1 2315 687 2315 687 1 ander_node_4
rlabel metal1 2168 687 2168 687 1 ander_node_3
rlabel metal1 2022 686 2022 686 1 ander_node_2
rlabel metal1 1886 685 1886 685 1 ander_node_1
rlabel metal2 2295 669 2295 669 1 A0
rlabel metal2 2149 669 2149 669 1 A1
rlabel metal2 2002 667 2002 667 1 A2
rlabel metal2 1874 662 1874 662 1 A3
rlabel metal1 2526 687 2526 687 1 ander_node_9
rlabel metal1 2660 687 2660 687 1 ander_node_10
rlabel metal1 2810 690 2810 690 1 ander_node_11
rlabel metal1 2954 687 2954 687 1 ander_node_12
rlabel metal1 2567 703 2567 703 1 A3_and_B3_nand
rlabel metal1 2695 704 2695 704 1 A2_and_B2_nand
rlabel metal1 2850 705 2850 705 1 A1_and_B1_nand
rlabel metal1 2990 705 2990 705 1 A0_and_B0_nand
rlabel metal1 2608 703 2608 703 1 A3_and_B3
rlabel metal1 2744 703 2744 703 1 A2_and_B2
rlabel metal1 2889 705 2889 705 1 A1_and_B1
rlabel metal1 3037 705 3037 705 1 A0_and_B0
rlabel metal1 1197 464 1197 464 1 compare_node_1
rlabel metal1 1058 464 1058 464 1 compare_node_2
rlabel metal1 912 465 912 465 1 compare_node_3
rlabel metal1 766 465 766 465 1 compare_node_4
rlabel metal1 757 359 757 359 1 compare_node_5
rlabel metal1 901 357 901 357 1 compare_node_6
rlabel metal1 1051 354 1051 354 1 compare_node_7
rlabel metal1 1194 354 1194 354 1 compare_node_8
rlabel metal1 1197 495 1197 495 1 compare_A3e_nand
rlabel metal1 1063 494 1063 494 1 compare_A2e_nand
rlabel metal1 917 493 917 493 1 compare_A1e_nand
rlabel metal1 769 497 769 497 1 compare_A0e_nand
rlabel metal1 761 390 761 390 1 compare_B0e_nand
rlabel metal1 906 387 906 387 1 compare_B1e_nand
rlabel metal1 1054 386 1054 386 1 compare_B2e_nand
rlabel metal1 1199 386 1199 386 1 compare_B3e_nand
rlabel metal1 1113 480 1113 480 1 compare_A3e
rlabel metal1 978 481 978 481 1 compare_A2e
rlabel metal1 834 481 834 481 1 compare_A1e
rlabel metal1 685 483 685 483 1 compare_A0e
rlabel metal1 677 375 677 375 1 compare_B0e
rlabel metal1 823 374 823 374 1 compare_B1e
rlabel metal1 972 371 972 371 1 compare_B2e
rlabel metal1 1117 372 1117 372 1 compare_B3e
rlabel pdiffusion 335 720 335 720 1 xnor_1
rlabel ndiffusion 335 680 335 680 1 xnor_2
rlabel metal1 396 709 396 709 1 xor_1
rlabel ndiffusion 417 720 417 720 1 xnor_3
rlabel pdiffusion 417 680 417 680 1 xnor_4
rlabel metal1 425 634 425 634 1 A3c
rlabel metal1 382 751 382 751 1 B3c
rlabel pdiffusion 330 498 330 498 1 xnor_5
rlabel ndiffusion 333 458 333 458 1 xnor_6
rlabel ndiffusion 416 498 416 498 1 xnor_7
rlabel pdiffusion 412 457 412 457 1 xnor_8
rlabel metal1 424 409 424 409 1 A2c
rlabel metal1 383 531 383 531 1 B2c
rlabel metal1 383 346 383 346 1 B1c
rlabel metal1 417 223 417 223 1 A1c
rlabel pdiffusion 335 312 335 312 1 xnor_9
rlabel ndiffusion 338 273 338 273 1 xnor_10
rlabel pdiffusion 416 273 416 273 1 xnor_11
rlabel ndiffusion 418 313 418 313 1 xnor_12
rlabel metal1 385 485 385 485 1 xor_2
rlabel metal1 390 301 390 301 1 xor_3
rlabel metal1 393 170 393 170 1 B0c
rlabel metal1 417 49 417 49 1 A0c
rlabel metal1 393 127 393 127 1 xor_4
rlabel pdiffusion 334 138 334 138 1 xnor_13
rlabel ndiffusion 336 97 336 97 1 xnor_14
rlabel ndiffusion 418 137 418 137 1 xnor_15
rlabel pdiffusion 418 98 418 98 1 xnor_16
rlabel ndiffusion 88 290 88 290 1 A_compare_B_node_3
rlabel ndiffusion 105 291 105 291 1 A_compare_B_node_2
rlabel ndiffusion 120 291 120 291 1 A_compare_B_node_1
rlabel metal1 5 315 5 315 3 A_equal_B
rlabel metal1 51 303 51 303 1 A_equal_B_c
rlabel metal1 94 373 94 373 1 A2e_xnor_B2e
rlabel metal1 223 711 223 711 1 A3e_xnor_B3e
rlabel metal1 222 303 222 303 1 A1e_xnor_B1e
rlabel metal1 223 127 223 127 1 A0e_xnor_B0e
rlabel metal2 2307 561 2307 561 1 B0
rlabel metal1 1214 712 1214 712 1 A_greater_B_node_1
rlabel metal1 1126 728 1126 728 1 A3_and_B3c
rlabel metal1 1211 744 1211 744 1 A3_nand_B3c
rlabel ndiffusion 1070 720 1070 720 1 A_greater_B_node_2
rlabel ndiffusion 1054 720 1054 720 1 A_greater_B_node_3
rlabel metal1 1024 728 1024 728 1 A3_eq_B3_A2_gt_B2_c
rlabel metal1 969 746 969 746 1 A3_eq_B3_A2_gt_B2
rlabel ndiffusion 928 721 928 721 1 A_greater_B_node_5
rlabel ndiffusion 907 722 907 722 1 A_greater_B_node_6
rlabel ndiffusion 891 720 891 720 1 A_greater_B_node_7
rlabel metal1 866 734 866 734 1 A3_eq_B3_A2_eq_B2_A1_gt_B1_c
rlabel metal1 812 747 812 747 1 A3_eq_B3_A2_eq_B2_A1_gt_B1
rlabel ndiffusion 734 723 734 723 1 A_greater_B_node_9
rlabel ndiffusion 715 722 715 722 1 A_greater_B_node_10
rlabel ndiffusion 699 722 699 722 1 A_greater_B_node_11
rlabel metal1 675 732 675 732 1 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0_c
rlabel metal1 622 746 622 746 1 A3_eq_B3_A2_eq_B2_A1_eq_B1_A0_gt_B0
rlabel ndiffusion 750 721 750 721 1 A_greater_B_node_8
rlabel pdiffusion 710 959 710 959 1 A_GT_B_node_1
rlabel pdiffusion 694 958 694 958 1 A_GT_B_node_2
rlabel pdiffusion 677 960 677 960 1 A_GT_B_node_3
rlabel metal1 750 933 750 933 1 A_GT_B_c
rlabel metal1 792 950 792 950 1 A_GT_B
rlabel metal1 948 1014 948 1014 1 A_LS_B_node_1
rlabel metal1 954 1045 954 1045 1 A_LS_B_nand
rlabel metal1 864 1031 864 1031 1 A_LS_B
rlabel metal1 2028 339 2028 339 1 D0_OR_D1_node
rlabel metal1 2027 365 2027 365 1 D0_OR_D1_node_2
rlabel metal1 2063 349 2063 349 1 D0_or_D1_c
rlabel metal1 2096 353 2096 353 1 D0_or_D1
rlabel metal1 2286 397 2286 397 1 adder_node1
rlabel metal1 2421 398 2421 398 1 adder_node2
rlabel metal1 2565 400 2565 400 1 adder_node3
rlabel metal1 2716 399 2716 399 1 adder_node4
rlabel metal1 2724 292 2724 292 1 adder_node5
rlabel metal1 2585 290 2585 290 1 adder_node6
rlabel metal1 2430 290 2430 290 1 adder_node7
rlabel metal1 2285 288 2285 288 1 adder_node8
rlabel metal1 2324 414 2324 414 1 Adder_A3ec
rlabel metal1 2463 413 2463 413 1 Adder_A2ec
rlabel metal1 2619 416 2619 416 1 Adder_A1ec
rlabel metal1 2754 415 2754 415 1 Adder_A0ec
rlabel metal1 2763 308 2763 308 1 Adder_B0ec
rlabel metal1 2635 307 2635 307 1 Adder_B1ec
rlabel metal1 2474 306 2474 306 1 Adder_B2ec
rlabel metal1 2325 306 2325 306 1 Adder_B3ec
rlabel metal1 2366 414 2366 414 1 adder_A3e
rlabel metal1 2502 413 2502 413 1 adder_A2e
rlabel metal1 2648 415 2648 415 1 adder_A1e
rlabel metal1 2795 415 2795 415 1 adder_A0e
rlabel metal1 2803 308 2803 308 1 adder_B0e
rlabel metal1 2661 307 2661 307 1 adder_B1e
rlabel metal1 2511 305 2511 305 1 adder_B2e
rlabel metal1 2367 306 2367 306 1 adder_B3e
rlabel metal1 2186 140 2186 140 1 B3ec_M
rlabel metal1 2186 -43 2186 -43 1 B2ec_M
rlabel metal1 2217 -216 2217 -216 1 B1ec_M
rlabel metal1 2235 -398 2235 -398 1 01ec_M
rlabel ndiffusion 2171 107 2171 107 1 adder_xor_node1
rlabel pdiffusion 2089 108 2089 108 1 adder_xor_node2
rlabel pdiffusion 2175 69 2175 69 1 adder_xor_node4
rlabel pdiffusion 2085 -75 2085 -75 1 adder_xor_node5
rlabel ndiffusion 2167 -75 2167 -75 1 adder_xor_node6
rlabel ndiffusion 2082 -113 2082 -113 1 adder_xor_node7
rlabel pdiffusion 2166 -114 2166 -114 1 adder_xor_node8
rlabel ndiffusion 2155 -249 2155 -249 1 adder_xor_node9
rlabel pdiffusion 2071 -249 2071 -249 1 adder_xor_node10
rlabel ndiffusion 2073 -285 2073 -285 1 adder_xor_node11
rlabel pdiffusion 2159 -288 2159 -288 1 adder_xor_node12
rlabel pdiffusion 2062 -432 2062 -432 1 adder_xor_node13
rlabel ndiffusion 2145 -431 2145 -431 1 adder_xor_node14
rlabel ndiffusion 2063 -471 2063 -471 1 adder_xor_node15
rlabel pdiffusion 2146 -472 2146 -472 1 adder_xor_node16
rlabel metal1 2119 96 2119 96 1 B3e_xor_M
rlabel metal1 2103 -99 2103 -99 1 B2e_xor_M
rlabel metal1 2090 -267 2090 -267 1 B1e_xor_M
rlabel metal1 2079 -454 2079 -454 1 B0e_xor_M
rlabel ndiffusion 2093 68 2093 68 1 adder_xor_node3
<< end >>
