magic
tech scmos
timestamp 1699167563
<< nwell >>
rect -50 1 34 31
<< ntransistor >>
rect -28 -22 -23 -17
rect -12 -22 -7 -17
rect 4 -22 9 -17
<< ptransistor >>
rect -28 14 -23 19
rect -12 14 -7 19
rect 4 14 9 19
<< ndiffusion >>
rect -31 -22 -28 -17
rect -23 -22 -20 -17
rect -15 -22 -12 -17
rect -7 -22 -4 -17
rect 1 -22 4 -17
rect 9 -22 12 -17
<< pdiffusion >>
rect -31 14 -28 19
rect -23 14 -12 19
rect -7 14 4 19
rect 9 14 12 19
<< ndcontact >>
rect -36 -22 -31 -17
rect -20 -22 -15 -17
rect -4 -22 1 -17
rect 12 -22 17 -17
<< pdcontact >>
rect -36 14 -31 19
rect 12 14 17 19
<< nsubstratencontact >>
rect 21 14 26 19
<< polysilicon >>
rect -28 19 -23 22
rect -12 19 -7 22
rect 4 19 9 22
rect -28 0 -23 14
rect -12 0 -7 14
rect 4 0 9 14
rect -27 -5 -23 0
rect -11 -5 -7 0
rect 5 -5 9 0
rect -28 -17 -23 -5
rect -12 -17 -7 -5
rect 4 -17 9 -5
rect -28 -25 -23 -22
rect -12 -25 -7 -22
rect 4 -25 9 -22
<< polycontact >>
rect -32 -5 -27 0
rect -16 -5 -11 0
rect 0 -5 5 0
<< metal1 >>
rect -50 30 34 35
rect -36 19 -31 30
rect 21 19 26 30
rect -35 -5 -32 0
rect -19 -5 -16 0
rect -3 -5 0 0
rect 12 -8 17 14
rect 37 5 52 9
rect 76 5 80 9
rect 37 -8 40 5
rect -20 -12 40 -8
rect -20 -17 -15 -12
rect 12 -17 17 -12
rect -36 -26 -31 -22
rect -4 -25 1 -22
rect 43 -25 48 -8
rect -4 -26 48 -25
rect -36 -29 48 -26
use not_without_labels  not_without_labels_0
timestamp 1699100137
transform 1 0 50 0 1 -1
box -16 -12 33 36
<< labels >>
rlabel metal1 -13 33 -13 33 5 Vdd!
rlabel metal1 -33 -4 -33 -4 1 input_A
rlabel metal1 -18 -3 -18 -3 1 input_B
rlabel metal1 -2 -3 -2 -3 1 input_C
rlabel metal1 15 -3 15 -3 1 v_output_nor_3
rlabel metal1 -15 -28 -15 -28 1 Gnd!
rlabel pdiffusion -1 17 -1 17 1 node_1
rlabel pdiffusion -18 17 -18 17 1 node_2
rlabel metal1 78 7 78 7 7 v_output_or_3
<< end >>
