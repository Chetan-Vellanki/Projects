.include "TSMC_180nm.txt"

* TESTING A 2:4 DECODER

.param supply_voltage = 1.5

.global Gnd
.global Vdd

VDD Vdd Gnd 'supply_voltage'
V_S0 S0 gnd PULSE(0 1.5 0 50p 50p 100n 200n)
V_S1 S1 gnd PULSE(0 1.5 0 50p 50p 50n 100n)

* SPICE3 file created from DECODER.ext - technology: scmos

.option scale=90n

M1000 DEC_D1_NAND S1c Vdd Vdd CMOSP w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1001 Vdd S0 DEC_D1_NAND Vdd CMOSP w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1002 DEC_D2_NAND S0c DEC_AND_NODE_3 Gnd CMOSN w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1003 Dec_AND_node_1 S1c Gnd Gnd CMOSN w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1004 DEC_AND_NODE_3 S1 Gnd Gnd CMOSN w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1005 S1c S1 Vdd Vdd CMOSP w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1006 S0c S0 Gnd Gnd CMOSN w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1007 D0 DEC_D0_NAND Gnd Gnd CMOSN w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1008 DEC_D3_NAND S1 Vdd Vdd CMOSP w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1009 D3 DEC_D3_NAND Vdd Vdd CMOSP w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1010 DEC_D1_NAND S1c Dec_AND_node_2 Gnd CMOSN w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1011 Dec_AND_node_2 S0 Gnd Gnd CMOSN w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1012 D1 DEC_D1_NAND Gnd Gnd CMOSN w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1013 D2 DEC_D2_NAND Gnd Gnd CMOSN w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1014 DEC_D3_NAND S1 DEC_AND_NODE_4 Gnd CMOSN w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
M1015 Vdd S0 DEC_D3_NAND Vdd CMOSP w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1016 D2 DEC_D2_NAND Vdd Vdd CMOSP w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1017 S0c S0 Vdd Vdd CMOSP w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1018 DEC_D0_NAND S0c Vdd Vdd CMOSP w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1019 D0 DEC_D0_NAND Vdd Vdd CMOSP w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1020 D1 DEC_D1_NAND Vdd Vdd CMOSP w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1021 DEC_AND_NODE_4 S0 Gnd Gnd CMOSN w=5 l=5
+  ad=35p pd=24u as=29.999998p ps=22u
M1022 S1c S1 Gnd Gnd CMOSN w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1023 DEC_D2_NAND S0c Vdd Vdd CMOSP w=5 l=5
+  ad=45p pd=23u as=35p ps=24u
M1024 D3 DEC_D3_NAND Gnd Gnd CMOSN w=5 l=5
+  ad=40p pd=26u as=35p ps=24u
M1025 Vdd S1 DEC_D2_NAND Vdd CMOSP w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1026 Vdd S1c DEC_D0_NAND Vdd CMOSP w=5 l=5
+  ad=35p pd=24u as=45p ps=23u
M1027 DEC_D0_NAND S0c Dec_AND_node_1 Gnd CMOSN w=5 l=5
+  ad=29.999998p pd=22u as=35p ps=24u
C0 DEC_D0_NAND Vdd 0.094023f
C1 Vdd Gnd 0.040225f
C2 DEC_D1_NAND Gnd 0.159401f
C3 D1 Gnd 0.051616f
C4 DEC_D0_NAND S1c 0.015311f
C5 DEC_D2_NAND DEC_AND_NODE_3 0.085282f
C6 S1 DEC_AND_NODE_4 0.088221f
C7 Vdd DEC_D1_NAND 0.094035f
C8 DEC_D2_NAND S0c 0.006448f
C9 D3 DEC_D3_NAND 0.030251f
C10 Gnd S1c 0.055406f
C11 S1 Gnd 0.142136f
C12 DEC_D1_NAND D1 0.030251f
C13 Vdd D1 0.04098f
C14 DEC_D0_NAND D0 0.030251f
C15 Vdd S1c 0.19269f
C16 S1 Vdd 0.201148f
C17 DEC_D1_NAND S1c 0.006448f
C18 Dec_AND_node_2 Gnd 0.077312f
C19 D0 Gnd 0.051616f
C20 DEC_D0_NAND Dec_AND_node_1 0.085282f
C21 DEC_AND_NODE_4 DEC_D3_NAND 0.085282f
C22 DEC_D0_NAND S0c 0.006448f
C23 Gnd DEC_D3_NAND 0.157853f
C24 Gnd DEC_AND_NODE_3 0.077196f
C25 S1 S1c 0.030251f
C26 DEC_AND_NODE_4 S0 0.089107f
C27 Dec_AND_node_1 Gnd 0.07683f
C28 DEC_D1_NAND Dec_AND_node_2 0.085282f
C29 Vdd D0 0.040884f
C30 DEC_D2_NAND D2 0.030251f
C31 Gnd S0 0.092334f
C32 Gnd S0c 0.051616f
C33 Vdd DEC_D3_NAND 0.094059f
C34 Dec_AND_node_2 S1c 0.088221f
C35 Vdd S0 0.202075f
C36 DEC_D1_NAND S0 0.015311f
C37 Vdd S0c 0.236061f
C38 S1 DEC_D3_NAND 0.006448f
C39 S1 DEC_AND_NODE_3 0.089107f
C40 Dec_AND_node_1 S1c 0.089107f
C41 S1c S0 0.07308f
C42 S1 S0 0.028532f
C43 S1c S0c 0.015985f
C44 S1 S0c 0.481731f
C45 Gnd DEC_D2_NAND 0.157853f
C46 Gnd D2 0.051616f
C47 D3 Gnd 0.051616f
C48 Vdd DEC_D2_NAND 0.094003f
C49 Dec_AND_node_2 S0 0.089107f
C50 Vdd D2 0.04098f
C51 Vdd D3 0.04098f
C52 DEC_D3_NAND S0 0.015311f
C53 DEC_AND_NODE_3 S0c 0.088221f
C54 DEC_D0_NAND Gnd 0.148342f
C55 Dec_AND_node_1 S0c 0.088221f
C56 S1 DEC_D2_NAND 0.015311f
C57 DEC_AND_NODE_4 Gnd 0.077062f
C58 S0 S0c 0.043542f
* C59 DEC_AND_NODE_4 0 0.248064f **FLOATING
* C60 D3 0 0.114466f **FLOATING
* C61 DEC_D3_NAND 0 0.516966f **FLOATING
* C62 DEC_AND_NODE_3 0 0.248064f **FLOATING
* C63 D2 0 0.114466f **FLOATING
* C64 DEC_D2_NAND 0 0.52029f **FLOATING
* C65 Dec_AND_node_2 0 0.248064f **FLOATING
* C66 S1 0 2.80331f **FLOATING
* C67 D1 0 0.104663f **FLOATING
* C68 DEC_D1_NAND 0 0.513722f **FLOATING
* C69 S0 0 7.95588f **FLOATING
* C70 Gnd 0 8.8184f **FLOATING
* C71 Dec_AND_node_1 0 0.248064f **FLOATING
* C72 D0 0 0.075352f **FLOATING
* C73 DEC_D0_NAND 0 0.520081f **FLOATING
* C74 S1c 0 4.39993f **FLOATING
* C75 S0c 0 5.11608f **FLOATING
* C76 Vdd 0 14.7872f **FLOATING


.tran 1n 1u

.control
run
plot v(S1)+10 v(S0)+8 v(D0)+6 v(D1)+4 v(D2)+2 v(D3)
.endc
.end