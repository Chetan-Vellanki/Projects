magic
tech scmos
timestamp 1701505937
<< nwell >>
rect 134 299 218 329
rect 225 309 271 328
rect 42 190 103 207
rect 117 174 163 193
rect 178 190 239 207
rect 253 174 299 193
rect 324 192 385 209
rect 399 176 445 195
rect -52 62 16 63
rect 235 62 247 64
rect 281 62 354 63
rect -106 43 16 62
rect 232 43 354 62
rect -37 36 16 43
rect 301 36 354 43
rect -36 35 16 36
rect 302 35 354 36
rect 46 24 61 29
rect 384 24 399 29
rect 46 15 98 24
rect 31 -4 98 15
rect 113 0 159 19
rect 384 15 436 24
rect 369 -4 436 15
rect 451 0 497 19
<< ntransistor >>
rect 251 294 256 299
rect 156 276 161 281
rect 172 276 177 281
rect 188 276 193 281
rect 62 167 67 172
rect 85 167 90 172
rect 198 167 203 172
rect 221 167 226 172
rect 344 169 349 174
rect 367 169 372 174
rect 143 159 148 164
rect 279 159 284 164
rect 425 161 430 166
rect 61 46 66 51
rect 79 46 84 51
rect 399 46 404 51
rect 417 46 422 51
rect -79 28 -74 33
rect 253 28 258 33
rect -22 7 -17 12
rect -4 7 1 12
rect 316 7 321 12
rect 334 7 339 12
rect 139 -15 144 -10
rect 477 -15 482 -10
<< ptransistor >>
rect 156 312 161 317
rect 172 312 177 317
rect 188 312 193 317
rect 251 316 256 321
rect 62 196 67 201
rect 85 196 90 201
rect 198 196 203 201
rect 221 196 226 201
rect 344 198 349 203
rect 367 198 372 203
rect 143 181 148 186
rect 279 181 284 186
rect 425 183 430 188
rect -79 50 -74 55
rect -22 46 -17 51
rect -4 46 1 51
rect 253 50 258 55
rect 316 46 321 51
rect 334 46 339 51
rect 61 7 66 12
rect 79 7 84 12
rect 139 7 144 12
rect 399 7 404 12
rect 417 7 422 12
rect 477 7 482 12
<< ndiffusion >>
rect 249 294 251 299
rect 256 294 259 299
rect 153 276 156 281
rect 161 276 164 281
rect 169 276 172 281
rect 177 276 180 281
rect 185 276 188 281
rect 193 276 196 281
rect 60 167 62 172
rect 67 167 69 172
rect 83 167 85 172
rect 90 167 92 172
rect 196 167 198 172
rect 203 167 205 172
rect 219 167 221 172
rect 226 167 228 172
rect 342 169 344 174
rect 349 169 351 174
rect 365 169 367 174
rect 372 169 374 174
rect 141 159 143 164
rect 148 159 151 164
rect 277 159 279 164
rect 284 159 287 164
rect 423 161 425 166
rect 430 161 433 166
rect 58 46 61 51
rect 66 46 79 51
rect 84 46 87 51
rect 396 46 399 51
rect 404 46 417 51
rect 422 46 425 51
rect -82 28 -79 33
rect -74 28 -72 33
rect 250 28 253 33
rect 258 28 260 33
rect -25 7 -22 12
rect -17 7 -4 12
rect 1 7 4 12
rect 313 7 316 12
rect 321 7 334 12
rect 339 7 342 12
rect 137 -15 139 -10
rect 144 -15 147 -10
rect 475 -15 477 -10
rect 482 -15 485 -10
<< pdiffusion >>
rect 153 312 156 317
rect 161 312 172 317
rect 177 312 188 317
rect 193 312 196 317
rect 249 316 251 321
rect 256 316 259 321
rect 60 196 62 201
rect 67 196 74 201
rect 79 196 85 201
rect 90 196 92 201
rect 196 196 198 201
rect 203 196 210 201
rect 215 196 221 201
rect 226 196 228 201
rect 342 198 344 203
rect 349 198 356 203
rect 361 198 367 203
rect 372 198 374 203
rect 141 181 143 186
rect 148 181 151 186
rect 277 181 279 186
rect 284 181 287 186
rect 423 183 425 188
rect 430 183 433 188
rect -82 50 -79 55
rect -74 50 -72 55
rect -25 46 -22 51
rect -17 46 -4 51
rect 1 46 4 51
rect 250 50 253 55
rect 258 50 260 55
rect 313 46 316 51
rect 321 46 334 51
rect 339 46 342 51
rect 58 7 61 12
rect 66 7 79 12
rect 84 7 87 12
rect 137 7 139 12
rect 144 7 147 12
rect 396 7 399 12
rect 404 7 417 12
rect 422 7 425 12
rect 475 7 477 12
rect 482 7 485 12
<< ndcontact >>
rect 244 294 249 299
rect 259 294 264 299
rect 148 276 153 281
rect 164 276 169 281
rect 180 276 185 281
rect 196 276 201 281
rect 55 167 60 172
rect 69 167 73 172
rect 79 167 83 172
rect 92 167 97 172
rect 191 167 196 172
rect 205 167 209 172
rect 215 167 219 172
rect 228 167 233 172
rect 337 169 342 174
rect 351 169 355 174
rect 361 169 365 174
rect 374 169 379 174
rect 136 159 141 164
rect 151 159 156 164
rect 272 159 277 164
rect 287 159 292 164
rect 418 161 423 166
rect 433 161 438 166
rect 53 46 58 51
rect 87 46 92 51
rect 391 46 396 51
rect 425 46 430 51
rect -87 28 -82 33
rect -72 28 -67 33
rect 245 28 250 33
rect 260 28 265 33
rect -30 7 -25 12
rect 4 7 9 12
rect 308 7 313 12
rect 342 7 347 12
rect 132 -15 137 -10
rect 147 -15 152 -10
rect 470 -15 475 -10
rect 485 -15 490 -10
<< pdcontact >>
rect 148 312 153 317
rect 196 312 201 317
rect 244 316 249 321
rect 259 316 264 321
rect 55 196 60 201
rect 74 196 79 201
rect 92 196 97 201
rect 191 196 196 201
rect 210 196 215 201
rect 228 196 233 201
rect 337 198 342 203
rect 356 198 361 203
rect 374 198 379 203
rect 136 181 141 186
rect 151 181 156 186
rect 272 181 277 186
rect 287 181 292 186
rect 418 183 423 188
rect 433 183 438 188
rect -87 50 -82 55
rect -72 50 -67 55
rect -30 46 -25 51
rect 4 46 9 51
rect 245 50 250 55
rect 260 50 265 55
rect 308 46 313 51
rect 342 46 347 51
rect 53 7 58 12
rect 87 7 92 12
rect 132 7 137 12
rect 147 7 152 12
rect 391 7 396 12
rect 425 7 430 12
rect 470 7 475 12
rect 485 7 490 12
<< nsubstratencontact >>
rect 205 312 210 317
rect 232 316 237 321
rect 46 196 51 201
rect 182 196 187 201
rect 328 198 333 203
rect 124 181 129 186
rect 260 181 265 186
rect 406 183 411 188
rect -60 50 -55 55
rect -42 46 -37 51
rect 272 50 277 55
rect 296 46 301 51
rect 38 5 43 10
rect 120 7 125 12
rect 376 5 381 10
rect 458 7 463 12
<< polysilicon >>
rect 251 321 256 324
rect 156 317 161 320
rect 172 317 177 320
rect 188 317 193 320
rect 156 281 161 312
rect 172 281 177 312
rect 188 281 193 312
rect 251 307 256 316
rect 252 303 256 307
rect 251 299 256 303
rect 251 289 256 294
rect 156 265 161 276
rect 172 265 177 276
rect 188 265 193 276
rect 62 201 67 215
rect 85 201 90 215
rect 198 201 203 215
rect 221 201 226 215
rect 344 203 349 217
rect 367 203 372 217
rect 62 172 67 196
rect 85 172 90 196
rect 143 186 148 189
rect 143 172 148 181
rect 198 172 203 196
rect 221 172 226 196
rect 279 186 284 189
rect 279 172 284 181
rect 344 174 349 198
rect 367 174 372 198
rect 425 188 430 191
rect 425 174 430 183
rect 144 168 148 172
rect 62 148 67 167
rect 85 148 90 167
rect 143 164 148 168
rect 280 168 284 172
rect 426 170 430 174
rect 143 154 148 159
rect 198 148 203 167
rect 221 148 226 167
rect 279 164 284 168
rect 279 154 284 159
rect 344 150 349 169
rect 367 150 372 169
rect 425 166 430 170
rect 425 156 430 161
rect -4 72 34 73
rect 39 72 84 73
rect -4 68 84 72
rect -79 55 -74 58
rect -22 51 -17 55
rect -4 51 1 68
rect 61 51 66 55
rect 79 51 84 68
rect 334 72 372 73
rect 377 72 422 73
rect 334 68 422 72
rect 253 55 258 58
rect -79 41 -74 50
rect 316 51 321 55
rect 334 51 339 68
rect 399 51 404 55
rect 417 51 422 68
rect -79 37 -75 41
rect -79 33 -74 37
rect -22 34 -17 46
rect -4 42 1 46
rect 61 34 66 46
rect 79 42 84 46
rect 253 41 258 50
rect 253 37 257 41
rect -21 29 1 34
rect 61 29 84 34
rect 253 33 258 37
rect 316 34 321 46
rect 334 42 339 46
rect 399 34 404 46
rect 417 42 422 46
rect -79 23 -74 28
rect -41 17 -17 22
rect -41 9 -36 17
rect -22 12 -17 17
rect -4 12 1 29
rect 61 12 66 16
rect 79 12 84 29
rect 317 29 339 34
rect 399 29 422 34
rect 253 23 258 28
rect 297 17 321 22
rect 139 12 144 15
rect -22 -11 -17 7
rect -4 1 1 7
rect 297 9 302 17
rect 316 12 321 17
rect 334 12 339 29
rect 399 12 404 16
rect 417 12 422 29
rect 477 12 482 15
rect 61 -11 66 7
rect -22 -16 66 -11
rect 79 -28 84 7
rect 139 -2 144 7
rect 140 -6 144 -2
rect 139 -10 144 -6
rect 316 -11 321 7
rect 334 1 339 7
rect 399 -11 404 7
rect 139 -20 144 -15
rect 316 -16 404 -11
rect 417 -28 422 7
rect 477 -2 482 7
rect 478 -6 482 -2
rect 477 -10 482 -6
rect 477 -20 482 -15
<< polycontact >>
rect 247 303 252 307
rect 156 258 161 265
rect 172 258 177 265
rect 188 258 193 265
rect 139 168 144 172
rect 62 142 67 148
rect 275 168 280 172
rect 421 170 426 174
rect 85 142 90 148
rect 198 142 203 148
rect 221 142 226 148
rect 344 144 349 150
rect 367 144 372 150
rect 34 72 39 77
rect 372 72 377 77
rect -75 37 -70 41
rect 257 37 262 41
rect -26 29 -21 34
rect 312 29 317 34
rect -41 4 -36 9
rect 297 4 302 9
rect 135 -6 140 -2
rect 79 -33 84 -28
rect 473 -6 478 -2
rect 417 -33 422 -28
<< metal1 >>
rect 131 328 273 333
rect -107 212 -102 213
rect 94 212 125 213
rect 131 212 137 328
rect 148 317 153 328
rect 205 317 210 328
rect 232 321 237 328
rect 244 321 249 328
rect 196 290 201 312
rect 259 307 264 316
rect 221 303 247 307
rect 259 303 310 307
rect 221 290 224 303
rect 259 299 264 303
rect 244 290 249 294
rect 164 286 224 290
rect 164 281 169 286
rect 196 281 201 286
rect 227 285 274 290
rect 148 273 153 276
rect 180 273 185 276
rect 227 273 232 285
rect 180 272 232 273
rect 153 269 232 272
rect 156 256 161 258
rect 172 256 177 258
rect 188 257 193 258
rect 376 214 404 215
rect 328 213 404 214
rect 230 212 404 213
rect -107 211 404 212
rect -107 209 379 211
rect -107 207 97 209
rect -107 206 52 207
rect -107 67 -102 206
rect 46 201 51 206
rect 55 201 60 207
rect 92 201 97 207
rect 117 208 233 209
rect 117 198 121 208
rect 182 207 233 208
rect 182 201 187 207
rect 74 186 79 196
rect 117 193 165 198
rect 191 201 196 207
rect 228 201 233 207
rect 253 198 257 209
rect 328 203 333 209
rect 337 203 342 209
rect 374 203 379 209
rect 399 200 403 211
rect 69 182 79 186
rect 124 186 129 193
rect 69 178 73 182
rect 136 186 141 193
rect 210 186 215 196
rect 253 193 301 198
rect 69 175 110 178
rect 69 172 73 175
rect 107 172 110 175
rect 151 172 156 181
rect 205 182 215 186
rect 260 186 265 193
rect 205 178 209 182
rect 272 186 277 193
rect 356 188 361 198
rect 399 196 473 200
rect 399 195 447 196
rect 205 175 246 178
rect 52 156 55 170
rect 97 167 99 170
rect 107 168 139 172
rect 151 168 168 172
rect 205 172 209 175
rect 243 172 246 175
rect 287 172 292 181
rect 351 184 361 188
rect 406 188 411 195
rect 351 180 355 184
rect 418 188 423 195
rect 351 177 392 180
rect 351 174 355 177
rect 389 174 392 177
rect 433 174 438 183
rect 79 164 82 167
rect 96 156 99 167
rect 151 164 156 168
rect 52 151 99 156
rect 136 155 141 159
rect 188 156 191 170
rect 233 167 235 170
rect 243 168 275 172
rect 287 168 309 172
rect 215 164 218 167
rect 232 156 235 167
rect 287 164 292 168
rect 131 150 166 155
rect 188 151 235 156
rect 62 141 67 142
rect 85 141 90 142
rect 162 129 166 150
rect 272 155 277 159
rect 334 158 337 172
rect 379 169 381 172
rect 389 170 421 174
rect 433 170 456 174
rect 361 166 364 169
rect 378 158 381 169
rect 433 166 438 170
rect 267 154 302 155
rect 267 150 315 154
rect 334 153 381 158
rect 418 157 423 161
rect 413 152 451 157
rect 296 149 315 150
rect 198 141 203 142
rect 221 141 226 142
rect 306 129 313 149
rect 344 143 349 144
rect 367 143 372 144
rect 442 132 451 152
rect 162 125 442 129
rect 162 124 452 125
rect -53 120 32 121
rect -53 117 85 120
rect 28 116 85 117
rect 85 105 90 115
rect 286 105 291 115
rect 442 105 443 110
rect 85 100 180 105
rect 34 79 171 84
rect 34 77 39 79
rect -107 63 11 67
rect -107 62 -52 63
rect -72 55 -67 62
rect -60 55 -55 62
rect -42 51 -37 63
rect -87 41 -82 50
rect -30 51 -25 63
rect 53 57 106 63
rect 53 51 58 57
rect -107 37 -82 41
rect -70 37 -52 41
rect -107 -27 -103 37
rect -87 33 -82 37
rect -47 34 -43 41
rect 4 40 9 46
rect 87 40 92 46
rect 4 35 21 40
rect 26 35 92 40
rect -47 29 -26 34
rect -72 24 -67 28
rect -97 19 -57 24
rect -62 -18 -57 19
rect 4 12 9 35
rect 53 29 56 32
rect 51 24 61 29
rect -41 1 -36 4
rect 53 12 58 24
rect -30 -18 -25 7
rect 87 12 92 35
rect 101 -18 106 57
rect 118 19 161 24
rect 120 12 125 19
rect 132 12 137 19
rect 147 -1 152 7
rect 166 -1 171 79
rect 132 -6 135 -2
rect 147 -6 171 -1
rect 147 -10 152 -6
rect -62 -19 106 -18
rect 132 -19 137 -15
rect -62 -23 155 -19
rect 101 -24 155 -23
rect -107 -32 62 -27
rect 21 -55 26 -40
rect 57 -37 62 -32
rect 79 -37 84 -33
rect 175 -31 180 100
rect 286 99 450 105
rect 286 83 291 99
rect 467 96 473 196
rect 493 111 498 165
rect 372 79 509 84
rect 372 77 377 79
rect 232 63 349 67
rect 232 62 281 63
rect 260 55 265 62
rect 272 55 277 62
rect 296 51 301 63
rect 245 41 250 50
rect 308 51 313 63
rect 391 57 444 63
rect 391 51 396 57
rect 124 -36 180 -31
rect 231 37 250 41
rect 262 37 286 41
rect 231 -27 235 37
rect 245 33 250 37
rect 291 34 295 41
rect 342 40 347 46
rect 342 35 360 40
rect 425 40 430 46
rect 366 35 430 40
rect 291 29 312 34
rect 260 24 265 28
rect 240 19 281 24
rect 276 -18 281 19
rect 342 12 347 35
rect 391 29 394 32
rect 389 24 399 29
rect 297 1 302 4
rect 391 12 396 24
rect 308 -18 313 7
rect 425 12 430 35
rect 439 -18 444 57
rect 456 19 499 24
rect 458 12 463 19
rect 470 12 475 19
rect 485 -1 490 7
rect 504 -1 509 79
rect 470 -6 473 -2
rect 485 -6 509 -1
rect 485 -10 490 -6
rect 281 -19 444 -18
rect 470 -19 475 -15
rect 281 -23 496 -19
rect 439 -24 496 -23
rect 231 -32 400 -27
rect 57 -42 84 -37
rect 179 -55 185 -52
rect 21 -58 185 -55
rect 360 -57 366 -41
rect 395 -37 400 -32
rect 417 -37 422 -33
rect 395 -42 422 -37
<< m2contact >>
rect 147 266 153 273
rect 156 251 161 256
rect 172 251 177 256
rect 188 252 193 257
rect 168 168 173 173
rect 77 159 82 164
rect 124 149 131 156
rect 309 168 314 173
rect 213 159 218 164
rect 62 134 67 141
rect 85 134 90 141
rect 260 149 267 156
rect 359 161 364 166
rect 456 169 461 174
rect 406 151 413 158
rect 198 134 203 141
rect 221 134 226 141
rect 344 136 349 143
rect 367 136 372 143
rect 442 125 454 132
rect -60 117 -53 124
rect 85 115 90 122
rect -2 108 5 113
rect 286 115 293 120
rect 443 105 452 112
rect 11 62 16 67
rect -52 36 -47 41
rect 21 35 26 40
rect 46 24 51 29
rect -41 -4 -36 1
rect 113 19 118 24
rect 127 -6 132 -1
rect 155 -24 162 -18
rect 21 -40 26 -35
rect 117 -36 124 -30
rect 493 105 502 111
rect 461 88 474 96
rect 286 75 293 83
rect 349 62 354 67
rect 286 36 291 41
rect 360 35 366 41
rect 384 24 389 29
rect 297 -4 302 1
rect 451 19 456 24
rect 465 -6 470 -1
rect 274 -24 281 -18
rect 496 -27 503 -18
rect 360 -41 366 -35
rect 178 -52 185 -44
<< metal2 >>
rect 107 273 153 274
rect 107 269 147 273
rect -60 124 -54 257
rect -2 113 5 258
rect 107 162 113 269
rect 156 239 161 251
rect 193 253 459 256
rect 172 247 177 251
rect 172 243 194 247
rect 156 234 173 239
rect 169 173 173 234
rect 190 232 194 243
rect 190 227 313 232
rect 309 173 313 227
rect 456 174 459 253
rect 82 159 113 162
rect 218 159 244 162
rect 364 161 390 164
rect 103 155 113 159
rect 103 150 124 155
rect 239 155 244 159
rect 385 157 390 161
rect 239 150 260 155
rect 385 152 406 157
rect 62 113 67 134
rect 85 122 90 134
rect 198 119 203 134
rect 90 115 203 119
rect 221 119 226 134
rect 221 115 286 119
rect 344 119 349 136
rect 293 115 349 119
rect -52 108 -2 113
rect 5 111 67 113
rect 367 111 372 136
rect 454 125 522 130
rect 5 108 372 111
rect -52 41 -47 108
rect 452 105 493 111
rect 19 88 461 96
rect 19 87 464 88
rect 19 67 24 87
rect 16 62 38 67
rect -41 -46 -36 -4
rect 21 -35 26 35
rect 32 29 38 62
rect 32 24 46 29
rect 113 24 118 87
rect 286 41 291 75
rect 357 67 362 87
rect 354 62 376 67
rect 38 10 43 24
rect 117 -6 127 -2
rect 117 -30 123 -6
rect 162 -24 274 -18
rect 117 -46 123 -36
rect -41 -51 123 -46
rect 297 -45 302 -4
rect 360 -35 366 35
rect 370 29 376 62
rect 370 24 384 29
rect 451 24 456 87
rect 376 10 381 24
rect 455 -6 465 -2
rect 185 -46 302 -45
rect 455 -46 461 -6
rect 517 -18 521 125
rect 503 -24 521 -18
rect 185 -50 461 -46
rect 297 -51 461 -50
<< end >>
